// This is the unpowered netlist.
module processor (Dataw_en,
    Serial_input,
    Serial_output,
    clk,
    hlt,
    reset,
    start,
    data_mem_addr,
    instr,
    instr_mem_addr,
    read_data,
    write_data);
 output Dataw_en;
 input Serial_input;
 output Serial_output;
 input clk;
 output hlt;
 input reset;
 input start;
 output [7:0] data_mem_addr;
 input [15:0] instr;
 output [12:0] instr_mem_addr;
 input [15:0] read_data;
 output [15:0] write_data;

 wire \Arithmetic_Logic_Unit.ALU_000.ALU_func[0] ;
 wire \Arithmetic_Logic_Unit.ALU_000.ALU_func[1] ;
 wire \Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i2 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[13].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[3].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.p_Z ;
 wire \Arithmetic_Logic_Unit.op ;
 wire \Control_unit1.instr_decoder1.A[0] ;
 wire \Control_unit1.instr_decoder1.A[1] ;
 wire \Control_unit1.instr_decoder1.A[2] ;
 wire \Control_unit1.instr_stage1[0] ;
 wire \Control_unit1.instr_stage1[10] ;
 wire \Control_unit1.instr_stage1[11] ;
 wire \Control_unit1.instr_stage1[12] ;
 wire \Control_unit1.instr_stage1[1] ;
 wire \Control_unit1.instr_stage1[2] ;
 wire \Control_unit1.instr_stage1[3] ;
 wire \Control_unit1.instr_stage1[4] ;
 wire \Control_unit1.instr_stage1[5] ;
 wire \Control_unit1.instr_stage1[6] ;
 wire \Control_unit1.instr_stage1[7] ;
 wire \Control_unit1.instr_stage1[8] ;
 wire \Control_unit1.instr_stage1[9] ;
 wire \Control_unit2.instr_decoder2.A[1] ;
 wire \Control_unit2.instr_decoder2.A[2] ;
 wire \Control_unit2.instr_stage2[10] ;
 wire \Control_unit2.instr_stage2[11] ;
 wire \Control_unit2.instr_stage2[12] ;
 wire \Control_unit2.instr_stage2[3] ;
 wire \Control_unit2.instr_stage2[4] ;
 wire \Control_unit2.instr_stage2[5] ;
 wire \Control_unit2.instr_stage2[6] ;
 wire \Control_unit2.instr_stage2[7] ;
 wire \Control_unit2.instr_stage2[8] ;
 wire \Control_unit2.instr_stage2[9] ;
 wire \Stack_pointer.SP[0] ;
 wire \Stack_pointer.SP[1] ;
 wire \Stack_pointer.SP[2] ;
 wire \Stack_pointer.SP[3] ;
 wire \Stack_pointer.SP[4] ;
 wire \Stack_pointer.SP[5] ;
 wire \Stack_pointer.SP[6] ;
 wire \Stack_pointer.SP[7] ;
 wire \Stack_pointer.SP_next[0] ;
 wire \Stack_pointer.SP_next[1] ;
 wire \Stack_pointer.SP_next[2] ;
 wire \Stack_pointer.SP_next[3] ;
 wire \Stack_pointer.SP_next[4] ;
 wire \Stack_pointer.SP_next[5] ;
 wire \Stack_pointer.SP_next[6] ;
 wire \Stack_pointer.SP_next[7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_opt_1_0_clk;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2382_ (.I(\Arithmetic_Logic_Unit.ALU_000.ALU_func[0] ),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2383_ (.I(_2078_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2384_ (.I(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2385_ (.I(\Arithmetic_Logic_Unit.ALU_000.ALU_func[1] ),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2386_ (.I(_2081_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2387_ (.I(_2082_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2388_ (.I(_2083_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2389_ (.I(\Control_unit2.instr_decoder2.A[2] ),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2390_ (.A1(\Arithmetic_Logic_Unit.op ),
    .A2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2391_ (.A1(_2080_),
    .A2(\Control_unit2.instr_decoder2.A[1] ),
    .A3(_2084_),
    .A4(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2392_ (.A1(_2079_),
    .A2(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2393_ (.I(\Control_unit2.instr_stage2[12] ),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2394_ (.A1(_2089_),
    .A2(\Control_unit2.instr_stage2[11] ),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2395_ (.A1(_2088_),
    .A2(_2090_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2396_ (.I(_2091_),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2397_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i3 ),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2398_ (.A1(\Arithmetic_Logic_Unit.ALU_000.ALU_func[0] ),
    .A2(\Arithmetic_Logic_Unit.ALU_000.ALU_func[1] ),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2399_ (.A1(_2080_),
    .A2(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2400_ (.I(_2094_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2401_ (.I(_2095_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2402_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i3 ),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2403_ (.A1(_2078_),
    .A2(_2081_),
    .B(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2404_ (.I(_2098_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2405_ (.A1(_2083_),
    .A2(_2097_),
    .B(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2406_ (.I(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2407_ (.I(_2081_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2408_ (.A1(_2101_),
    .A2(_2102_),
    .B(_2093_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2409_ (.I(_2103_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2410_ (.A1(_2092_),
    .A2(_2096_),
    .A3(_2100_),
    .A4(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2411_ (.I(_2092_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2412_ (.I(_2094_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2413_ (.I(_2107_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2414_ (.I0(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ),
    .I1(_2078_),
    .S(_2081_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2415_ (.I(_2109_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2416_ (.A1(_2092_),
    .A2(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2417_ (.A1(_2106_),
    .A2(_2108_),
    .B1(_2100_),
    .B2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2418_ (.A1(_2105_),
    .A2(_2112_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2419_ (.I(\Control_unit1.instr_decoder1.A[0] ),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2420_ (.A1(\Control_unit1.instr_decoder1.A[2] ),
    .A2(\Control_unit1.instr_decoder1.A[1] ),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2421_ (.A1(\Control_unit1.instr_stage1[3] ),
    .A2(\Control_unit1.instr_stage1[1] ),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2422_ (.A1(_2114_),
    .A2(\Control_unit1.instr_stage1[2] ),
    .A3(_2115_),
    .A4(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2423_ (.I0(net37),
    .I1(net1),
    .S(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2424_ (.I(_2079_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2425_ (.A1(_2083_),
    .A2(_2118_),
    .B(_2119_),
    .C(_2101_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2426_ (.I(net37),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2427_ (.I(net1),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2428_ (.I0(_2121_),
    .I1(_2122_),
    .S(_2117_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2429_ (.I(_2102_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2430_ (.A1(_2078_),
    .A2(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2431_ (.I(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2432_ (.A1(_2079_),
    .A2(_2123_),
    .B(_2126_),
    .C(_2080_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2433_ (.A1(_2120_),
    .A2(_2127_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2434_ (.A1(_2113_),
    .A2(_2128_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2435_ (.I(_2102_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2436_ (.I(_2130_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2437_ (.I(_2131_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2438_ (.I(_2132_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2439_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2440_ (.I(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2441_ (.I(_2093_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2442_ (.I(_2136_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2443_ (.I(_2125_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2444_ (.I(_2138_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2445_ (.A1(_2133_),
    .A2(_2106_),
    .B1(_2135_),
    .B2(_2137_),
    .C1(_2139_),
    .C2(_2118_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2446_ (.I(\Arithmetic_Logic_Unit.op ),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2447_ (.I(_2141_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2448_ (.I(_2142_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2449_ (.I0(_2129_),
    .I1(_2140_),
    .S(_2143_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2450_ (.I(_2144_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2451_ (.I(_2145_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2452_ (.I(_2146_),
    .ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2453_ (.I(_2141_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2454_ (.I(_2147_),
    .Z(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2455_ (.I(_2095_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2456_ (.I(_2103_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2457_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2458_ (.I(_2098_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2459_ (.A1(_2082_),
    .A2(_2151_),
    .B(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _2460_ (.A1(_2134_),
    .A2(_2149_),
    .A3(_2150_),
    .A4(_2153_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2461_ (.I(_2109_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2462_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ),
    .A2(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2463_ (.A1(_2134_),
    .A2(_2096_),
    .B1(_2156_),
    .B2(_2153_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2464_ (.A1(_2154_),
    .A2(_2157_),
    .Z(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2465_ (.I(_2112_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2466_ (.A1(_2159_),
    .A2(_2128_),
    .B(_2105_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2467_ (.A1(_2158_),
    .A2(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2468_ (.I(_2142_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2469_ (.I(_2132_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2470_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2471_ (.I(_2164_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2472_ (.I(_2136_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(_2166_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2474_ (.A1(_2163_),
    .A2(_2135_),
    .B1(_2165_),
    .B2(_2167_),
    .C1(_2139_),
    .C2(_2106_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2475_ (.A1(_2162_),
    .A2(_2168_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2476_ (.A1(_2148_),
    .A2(_2161_),
    .B(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2477_ (.I(_2170_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2478_ (.I(_2171_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2479_ (.I(_2172_),
    .ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2480_ (.A1(_2113_),
    .A2(_2158_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2481_ (.A1(_2092_),
    .A2(_2096_),
    .A3(_2100_),
    .A4(_2104_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2482_ (.A1(_2174_),
    .A2(_2154_),
    .A3(_2157_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2483_ (.A1(_2128_),
    .A2(_2173_),
    .B(_2175_),
    .C(_2154_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2484_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2485_ (.A1(_2082_),
    .A2(_2177_),
    .B(_2099_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2486_ (.A1(_2164_),
    .A2(_2149_),
    .A3(_2150_),
    .A4(_2178_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2487_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ),
    .A2(_2110_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2488_ (.A1(_2164_),
    .A2(_2096_),
    .B1(_2180_),
    .B2(_2178_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2489_ (.A1(_2179_),
    .A2(_2181_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2490_ (.A1(_2176_),
    .A2(_2182_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2491_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[3].i3 ),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2492_ (.I(_2184_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2493_ (.A1(_2163_),
    .A2(_2165_),
    .B1(_2185_),
    .B2(_2167_),
    .C1(_2139_),
    .C2(_2135_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(_2162_),
    .A2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2495_ (.A1(_2148_),
    .A2(_2183_),
    .B(_2187_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2496_ (.I(_2188_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2497_ (.I(_2189_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2498_ (.I(_2190_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2499_ (.I(_2107_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2500_ (.A1(_2184_),
    .A2(_2110_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2501_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[3].i3 ),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2502_ (.A1(_2082_),
    .A2(_2193_),
    .B(_2098_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2503_ (.A1(_2184_),
    .A2(_2191_),
    .B1(_2192_),
    .B2(_2194_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2504_ (.A1(_2184_),
    .A2(_2107_),
    .A3(_2150_),
    .A4(_2194_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2505_ (.I(_2196_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2506_ (.A1(_2195_),
    .A2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(_2128_),
    .A2(_2173_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2508_ (.A1(_2134_),
    .A2(_2191_),
    .A3(_2104_),
    .A4(_2153_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2509_ (.A1(_2200_),
    .A2(_2179_),
    .A3(_2181_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2510_ (.A1(_2175_),
    .A2(_2179_),
    .A3(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2511_ (.A1(_2199_),
    .A2(_2182_),
    .B(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2512_ (.A1(_2198_),
    .A2(_2203_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2513_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2514_ (.I(_2205_),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2515_ (.I(_2166_),
    .Z(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2516_ (.I(_2138_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2517_ (.A1(_2163_),
    .A2(_2185_),
    .B1(_2206_),
    .B2(_2207_),
    .C1(_2208_),
    .C2(_2165_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2518_ (.I0(_2204_),
    .I1(_2209_),
    .S(_2162_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2519_ (.I(_2210_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2520_ (.I(_2211_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2521_ (.I(_2212_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2522_ (.A1(_2154_),
    .A2(_2157_),
    .A3(_2179_),
    .A4(_2181_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2523_ (.A1(_2105_),
    .A2(_2112_),
    .A3(_2195_),
    .A4(_2197_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2524_ (.A1(_2120_),
    .A2(_2127_),
    .A3(_2213_),
    .A4(_2214_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2525_ (.A1(_2164_),
    .A2(_2108_),
    .A3(_2104_),
    .A4(_2178_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2526_ (.A1(_2216_),
    .A2(_2195_),
    .A3(_2196_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2527_ (.A1(_2175_),
    .A2(_2197_),
    .A3(_2201_),
    .A4(_2217_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2528_ (.A1(_2205_),
    .A2(_2149_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2529_ (.A1(_2130_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2530_ (.A1(_2205_),
    .A2(_2155_),
    .B1(_2220_),
    .B2(_2099_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2531_ (.A1(_2219_),
    .A2(_2221_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2532_ (.I(_2222_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2533_ (.A1(_2215_),
    .A2(_2218_),
    .B(_2223_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2534_ (.A1(_2120_),
    .A2(_2127_),
    .A3(_2213_),
    .A4(_2214_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2535_ (.A1(_2175_),
    .A2(_2197_),
    .A3(_2201_),
    .A4(_2217_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2536_ (.A1(_2225_),
    .A2(_2226_),
    .A3(_2222_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2537_ (.A1(_2224_),
    .A2(_2227_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2538_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2539_ (.A1(_2229_),
    .A2(_2166_),
    .B1(_2138_),
    .B2(_2185_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2540_ (.A1(_2142_),
    .A2(_2220_),
    .A3(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2541_ (.A1(_2147_),
    .A2(_2228_),
    .B(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2542_ (.I(_2232_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2543_ (.I(_2162_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2544_ (.I(_2107_),
    .Z(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2545_ (.A1(_2205_),
    .A2(_2234_),
    .A3(_2221_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2546_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ),
    .A2(_2095_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2547_ (.A1(_2130_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2548_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ),
    .A2(_2109_),
    .B1(_2237_),
    .B2(_2152_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2549_ (.A1(_2236_),
    .A2(_2238_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2550_ (.I(_2239_),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2551_ (.A1(_2235_),
    .A2(_2224_),
    .A3(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2552_ (.A1(_2222_),
    .A2(_2239_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2553_ (.A1(_2225_),
    .A2(_2226_),
    .B(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2554_ (.A1(_2235_),
    .A2(_2240_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2555_ (.I(_2244_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2556_ (.A1(_2243_),
    .A2(_2245_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2557_ (.A1(_2241_),
    .A2(_2246_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2558_ (.I(_2143_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2559_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2560_ (.I(_2249_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2561_ (.I(_2137_),
    .Z(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2562_ (.I(_2125_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2563_ (.I(_2252_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2564_ (.A1(_2250_),
    .A2(_2251_),
    .B1(_2253_),
    .B2(_2206_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2565_ (.A1(_2248_),
    .A2(_2237_),
    .A3(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2566_ (.A1(_2233_),
    .A2(_2247_),
    .B(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2567_ (.I(_2256_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2568_ (.I(_2257_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2569_ (.I(_2143_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2570_ (.I(_2191_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2571_ (.I(_2259_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2572_ (.I(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2573_ (.A1(_2229_),
    .A2(_2261_),
    .A3(_2238_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2574_ (.A1(_2249_),
    .A2(_2095_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2575_ (.A1(_2130_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2576_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ),
    .A2(_2155_),
    .B1(_2264_),
    .B2(_2152_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2577_ (.A1(_2263_),
    .A2(_2265_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2578_ (.I(_2266_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2579_ (.I(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2580_ (.A1(_2262_),
    .A2(_2243_),
    .A3(_2245_),
    .A4(_2268_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2581_ (.A1(_2262_),
    .A2(_2243_),
    .A3(_2245_),
    .B(_2268_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2582_ (.A1(_2269_),
    .A2(_2270_),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2583_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2584_ (.I(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2585_ (.I(_2229_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2586_ (.A1(_2273_),
    .A2(_2251_),
    .B1(_2253_),
    .B2(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2587_ (.A1(_2148_),
    .A2(_2264_),
    .A3(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2588_ (.A1(_2258_),
    .A2(_2271_),
    .B(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2589_ (.I(_2277_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2590_ (.I(_2278_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2591_ (.I(_2147_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2592_ (.I(_2279_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2593_ (.A1(_2124_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2594_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2595_ (.I(_2282_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2596_ (.A1(_2283_),
    .A2(_2167_),
    .B1(_2208_),
    .B2(_2249_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2597_ (.A1(_2281_),
    .A2(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2598_ (.A1(_2272_),
    .A2(_2149_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2599_ (.A1(_2272_),
    .A2(_2110_),
    .B1(_2281_),
    .B2(_2099_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2600_ (.A1(_2286_),
    .A2(_2287_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2601_ (.A1(_2249_),
    .A2(_2259_),
    .A3(_2265_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2602_ (.I(_2289_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2603_ (.A1(_2229_),
    .A2(_2234_),
    .A3(_2238_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2604_ (.A1(_2291_),
    .A2(_2267_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2605_ (.A1(_2245_),
    .A2(_2290_),
    .A3(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2606_ (.A1(_2224_),
    .A2(_2240_),
    .A3(_2267_),
    .B(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2607_ (.A1(_2288_),
    .A2(_2294_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2608_ (.A1(_2280_),
    .A2(_2295_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2609_ (.A1(_2280_),
    .A2(_2285_),
    .B(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2610_ (.I(_2297_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2611_ (.I(_2298_),
    .ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2612_ (.A1(_2222_),
    .A2(_2240_),
    .A3(_2267_),
    .A4(_2288_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2613_ (.A1(_2215_),
    .A2(_2218_),
    .B(_2299_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2614_ (.A1(_2272_),
    .A2(_2259_),
    .A3(_2287_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2615_ (.A1(_2289_),
    .A2(_2288_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2616_ (.A1(_2244_),
    .A2(_2301_),
    .A3(_2292_),
    .A4(_2302_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2617_ (.A1(_2282_),
    .A2(_2234_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2618_ (.I(_2155_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2619_ (.A1(_2131_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2620_ (.I(_2152_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2621_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ),
    .A2(_2305_),
    .B1(_2306_),
    .B2(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2622_ (.A1(_2304_),
    .A2(_2308_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2623_ (.A1(_2300_),
    .A2(_2303_),
    .B(_2309_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2624_ (.A1(_2266_),
    .A2(_2288_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2625_ (.A1(_2225_),
    .A2(_2226_),
    .B(_2242_),
    .C(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _2626_ (.A1(_2244_),
    .A2(_2301_),
    .A3(_2292_),
    .A4(_2302_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2627_ (.A1(_2304_),
    .A2(_2308_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2628_ (.A1(_2312_),
    .A2(_2313_),
    .A3(_2314_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2629_ (.A1(_2310_),
    .A2(_2315_),
    .B(_2280_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2630_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2631_ (.I(_2317_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2632_ (.A1(_2133_),
    .A2(_2283_),
    .B1(_2318_),
    .B2(_2137_),
    .C1(_2252_),
    .C2(_2273_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2633_ (.A1(_2258_),
    .A2(_2319_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2634_ (.A1(_2316_),
    .A2(_2320_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2635_ (.I(_2321_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2636_ (.I(_2322_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2637_ (.A1(_2282_),
    .A2(_2259_),
    .A3(_2308_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2638_ (.A1(_2317_),
    .A2(_2191_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(_2124_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2640_ (.A1(_2317_),
    .A2(_2305_),
    .B1(_2325_),
    .B2(_2307_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2641_ (.A1(_2324_),
    .A2(_2326_),
    .Z(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2642_ (.A1(_2323_),
    .A2(_2327_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2643_ (.A1(_2309_),
    .A2(_2327_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2644_ (.A1(_2312_),
    .A2(_2313_),
    .B(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2645_ (.A1(_2323_),
    .A2(_2327_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2646_ (.A1(_2310_),
    .A2(_2328_),
    .B(_2330_),
    .C(_2331_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2647_ (.A1(_2133_),
    .A2(_2318_),
    .B1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ),
    .B2(_2166_),
    .C1(_2252_),
    .C2(_2282_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2648_ (.I0(_2332_),
    .I1(_2333_),
    .S(_2143_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2649_ (.I(_2334_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2650_ (.I(_2335_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2651_ (.I(_2336_),
    .ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2652_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ),
    .Z(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2653_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2654_ (.A1(_2083_),
    .A2(_2338_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2655_ (.A1(_2337_),
    .A2(_2137_),
    .B1(_2252_),
    .B2(_2318_),
    .C(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2656_ (.A1(_2248_),
    .A2(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2657_ (.I(_2234_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2658_ (.A1(_2317_),
    .A2(_2342_),
    .A3(_2326_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2659_ (.A1(_2343_),
    .A2(_2331_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2660_ (.I(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2661_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ),
    .A2(_2108_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2662_ (.A1(_2101_),
    .A2(_2136_),
    .A3(_2339_),
    .B1(_2150_),
    .B2(_2338_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2663_ (.A1(_2346_),
    .A2(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2664_ (.A1(_2330_),
    .A2(_2345_),
    .B(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2665_ (.A1(_2300_),
    .A2(_2303_),
    .B(_2309_),
    .C(_2327_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2666_ (.I(_2348_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2667_ (.A1(_2350_),
    .A2(_2351_),
    .A3(_2344_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2668_ (.A1(_2349_),
    .A2(_2352_),
    .B(_2280_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2669_ (.A1(_2341_),
    .A2(_2353_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2670_ (.I(_2354_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2671_ (.I(_2355_),
    .ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2672_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ),
    .A2(_2108_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2673_ (.A1(_2124_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2674_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ),
    .A2(_2305_),
    .B1(_2357_),
    .B2(_2307_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2675_ (.A1(_2356_),
    .A2(_2358_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2676_ (.A1(_2346_),
    .A2(_2347_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2677_ (.A1(_2343_),
    .A2(_2348_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2678_ (.A1(_2331_),
    .A2(_2360_),
    .A3(_2361_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2679_ (.A1(_2350_),
    .A2(_2351_),
    .B(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2680_ (.A1(_2359_),
    .A2(_2363_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2681_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2682_ (.I(_2365_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2683_ (.I(_2357_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2684_ (.A1(_2366_),
    .A2(_2136_),
    .B1(_2138_),
    .B2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ),
    .C(_2367_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2685_ (.A1(_2142_),
    .A2(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2686_ (.A1(_2147_),
    .A2(_2364_),
    .B(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2687_ (.I(_2370_),
    .ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2688_ (.A1(_2365_),
    .A2(_2342_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2689_ (.I(_2305_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2690_ (.A1(_2131_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2691_ (.I(_2307_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2692_ (.A1(_2365_),
    .A2(_2372_),
    .B1(_2373_),
    .B2(_2374_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2693_ (.A1(_2371_),
    .A2(_2375_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2694_ (.I(_2376_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2695_ (.A1(_2348_),
    .A2(_2359_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2696_ (.A1(_2329_),
    .A2(_2378_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2697_ (.A1(_2300_),
    .A2(_2303_),
    .B(_2379_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2698_ (.A1(_2337_),
    .A2(_2260_),
    .A3(_2358_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2699_ (.A1(_2360_),
    .A2(_2359_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2700_ (.A1(_2331_),
    .A2(_2381_),
    .A3(_2361_),
    .A4(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2701_ (.A1(_2377_),
    .A2(_2380_),
    .A3(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2702_ (.A1(_2312_),
    .A2(_2313_),
    .B(_2329_),
    .C(_2378_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2703_ (.I(_0560_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2704_ (.A1(_0562_),
    .A2(_0563_),
    .B(_2376_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2705_ (.A1(_0561_),
    .A2(_0564_),
    .B(_2279_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2706_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[13].i3 ),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2707_ (.I(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2708_ (.A1(_2163_),
    .A2(_2366_),
    .B1(_0567_),
    .B2(_2167_),
    .C1(_2139_),
    .C2(_2337_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2709_ (.A1(_2148_),
    .A2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2710_ (.A1(_0565_),
    .A2(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2711_ (.I(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2712_ (.I(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2713_ (.I(_0572_),
    .ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2714_ (.A1(_2380_),
    .A2(_0560_),
    .B(_2377_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2715_ (.A1(_2365_),
    .A2(_2261_),
    .A3(_2375_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2716_ (.A1(_2131_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[13].i3 ),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2717_ (.A1(_0566_),
    .A2(_2372_),
    .B1(_0575_),
    .B2(_2374_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2718_ (.A1(_0566_),
    .A2(_2342_),
    .A3(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2719_ (.I(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2720_ (.A1(_0566_),
    .A2(_2342_),
    .B(_0576_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2721_ (.A1(_0578_),
    .A2(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2722_ (.A1(_0574_),
    .A2(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2723_ (.A1(_2376_),
    .A2(_0580_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2724_ (.A1(_0562_),
    .A2(_0563_),
    .B(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2725_ (.A1(_0574_),
    .A2(_0580_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2726_ (.A1(_0573_),
    .A2(_0581_),
    .B(_0583_),
    .C(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2727_ (.I(_2133_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2728_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2729_ (.I(_0587_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2730_ (.A1(_0586_),
    .A2(_0567_),
    .B1(_0588_),
    .B2(_2207_),
    .C1(_2208_),
    .C2(_2366_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2731_ (.A1(_2258_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2732_ (.A1(_2258_),
    .A2(_0585_),
    .B(_0590_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2733_ (.I(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2734_ (.I(_0592_),
    .ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2735_ (.A1(_2132_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2736_ (.A1(_0587_),
    .A2(_2372_),
    .B1(_0593_),
    .B2(_2374_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2737_ (.A1(_0587_),
    .A2(_2260_),
    .A3(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2738_ (.I(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2739_ (.A1(_0587_),
    .A2(_2260_),
    .B(_0594_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2740_ (.A1(_0596_),
    .A2(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2741_ (.A1(_0578_),
    .A2(_0583_),
    .A3(_0584_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2742_ (.A1(_0598_),
    .A2(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2743_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i2 ),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2744_ (.A1(_0586_),
    .A2(_0588_),
    .B1(_0601_),
    .B2(_2207_),
    .C1(_2208_),
    .C2(_0567_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2745_ (.I0(_0600_),
    .I1(_0602_),
    .S(_2248_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2746_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2747_ (.I(_0604_),
    .ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2748_ (.A1(_0577_),
    .A2(_0598_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2749_ (.A1(_0562_),
    .A2(_0563_),
    .B(_0582_),
    .C(_0598_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2750_ (.A1(_0584_),
    .A2(_0596_),
    .A3(_0605_),
    .A4(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2751_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i2 ),
    .A2(_2261_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2752_ (.A1(_2132_),
    .A2(_0601_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2753_ (.A1(_0601_),
    .A2(_2372_),
    .B1(_0609_),
    .B2(_2374_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2754_ (.A1(_0607_),
    .A2(_0608_),
    .A3(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2755_ (.I(_0601_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2756_ (.A1(_0586_),
    .A2(_0612_),
    .B1(_2207_),
    .B2(_2118_),
    .C1(_2253_),
    .C2(_0588_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2757_ (.I0(_0611_),
    .I1(_0613_),
    .S(_2248_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2758_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2759_ (.I(_0615_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2760_ (.I(\Control_unit2.instr_decoder2.A[1] ),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2761_ (.A1(_2141_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.p_Z ),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2762_ (.A1(\Control_unit2.instr_decoder2.A[2] ),
    .A2(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2763_ (.A1(_0616_),
    .A2(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2764_ (.I(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2765_ (.I(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2766_ (.I(_0620_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2767_ (.A1(\Control_unit1.instr_decoder1.A[0] ),
    .A2(\Control_unit1.instr_stage1[2] ),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2768_ (.A1(\Control_unit1.instr_stage1[1] ),
    .A2(_2115_),
    .A3(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2769_ (.A1(\Control_unit1.instr_stage1[0] ),
    .A2(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2770_ (.A1(\Control_unit1.instr_stage1[12] ),
    .A2(\Control_unit1.instr_stage1[11] ),
    .A3(_0625_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2771_ (.A1(\Control_unit1.instr_decoder1.A[2] ),
    .A2(\Control_unit1.instr_decoder1.A[1] ),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2772_ (.A1(_0626_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2773_ (.A1(\Stack_pointer.SP[0] ),
    .A2(_0622_),
    .A3(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2774_ (.I(_0626_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2775_ (.I(_0627_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2776_ (.I(_0619_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2777_ (.A1(\Stack_pointer.SP[0] ),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2778_ (.A1(\Control_unit1.instr_stage1[3] ),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2779_ (.A1(\Stack_pointer.SP[0] ),
    .A2(_0621_),
    .B(_0629_),
    .C(_0634_),
    .ZN(\Stack_pointer.SP_next[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2780_ (.I(_0628_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2781_ (.A1(\Stack_pointer.SP[1] ),
    .A2(_0621_),
    .A3(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2782_ (.I(_0626_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2783_ (.I(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2784_ (.I(_0627_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2785_ (.I(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2786_ (.A1(\Stack_pointer.SP[1] ),
    .A2(_0622_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2787_ (.I(_0620_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2788_ (.A1(\Stack_pointer.SP[1] ),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2789_ (.A1(\Control_unit1.instr_stage1[4] ),
    .A2(_0638_),
    .B1(_0640_),
    .B2(_0641_),
    .C(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2790_ (.A1(_0636_),
    .A2(_0644_),
    .ZN(\Stack_pointer.SP_next[1] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2791_ (.A1(\Stack_pointer.SP[2] ),
    .A2(_0621_),
    .A3(_0635_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2792_ (.A1(\Stack_pointer.SP[2] ),
    .A2(_0622_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2793_ (.A1(\Stack_pointer.SP[2] ),
    .A2(_0642_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2794_ (.A1(\Control_unit1.instr_stage1[5] ),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0646_),
    .C(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2795_ (.A1(_0645_),
    .A2(_0648_),
    .ZN(\Stack_pointer.SP_next[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2796_ (.A1(\Stack_pointer.SP[3] ),
    .A2(_0621_),
    .A3(_0635_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2797_ (.A1(\Stack_pointer.SP[3] ),
    .A2(_0642_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2798_ (.I(_0619_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2799_ (.A1(\Stack_pointer.SP[3] ),
    .A2(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2800_ (.A1(\Control_unit1.instr_stage1[6] ),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0650_),
    .C(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2801_ (.A1(_0649_),
    .A2(_0653_),
    .ZN(\Stack_pointer.SP_next[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2802_ (.A1(\Stack_pointer.SP[4] ),
    .A2(_0622_),
    .A3(_0635_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2803_ (.A1(\Stack_pointer.SP[4] ),
    .A2(_0642_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2804_ (.A1(\Stack_pointer.SP[4] ),
    .A2(_0651_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2805_ (.A1(\Control_unit1.instr_stage1[7] ),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0655_),
    .C(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2806_ (.A1(_0654_),
    .A2(_0657_),
    .ZN(\Stack_pointer.SP_next[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2807_ (.A1(\Stack_pointer.SP[5] ),
    .A2(_0632_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2808_ (.A1(\Stack_pointer.SP[5] ),
    .A2(_0651_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2809_ (.A1(\Control_unit1.instr_stage1[8] ),
    .A2(_0637_),
    .B1(_0639_),
    .B2(_0658_),
    .C(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2810_ (.A1(_0638_),
    .A2(_0640_),
    .A3(_0658_),
    .B(_0660_),
    .ZN(\Stack_pointer.SP_next[5] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2811_ (.A1(\Stack_pointer.SP[6] ),
    .A2(_0632_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2812_ (.A1(\Stack_pointer.SP[6] ),
    .A2(_0651_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2813_ (.A1(\Control_unit1.instr_stage1[9] ),
    .A2(_0637_),
    .B1(_0639_),
    .B2(_0661_),
    .C(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2814_ (.A1(_0638_),
    .A2(_0640_),
    .A3(_0661_),
    .B(_0663_),
    .ZN(\Stack_pointer.SP_next[6] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2815_ (.A1(\Stack_pointer.SP[7] ),
    .A2(_0620_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2816_ (.A1(\Stack_pointer.SP[7] ),
    .A2(_0632_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2817_ (.A1(\Control_unit1.instr_stage1[10] ),
    .A2(_0637_),
    .B1(_0639_),
    .B2(_0664_),
    .C(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2818_ (.A1(_0638_),
    .A2(_0640_),
    .A3(_0664_),
    .B(_0666_),
    .ZN(\Stack_pointer.SP_next[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2819_ (.I(_0618_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2820_ (.A1(_2086_),
    .A2(_0667_),
    .B(_0616_),
    .ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2821_ (.I(\Control_unit1.instr_decoder1.A[2] ),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2822_ (.A1(_0668_),
    .A2(\Control_unit1.instr_decoder1.A[1] ),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2823_ (.A1(\Control_unit1.instr_decoder1.A[0] ),
    .A2(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2824_ (.I(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2825_ (.I(\Stack_pointer.SP[0] ),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2826_ (.A1(\Control_unit1.instr_stage1[12] ),
    .A2(\Control_unit1.instr_stage1[11] ),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2827_ (.A1(_0625_),
    .A2(_0673_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2828_ (.A1(_0672_),
    .A2(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2829_ (.A1(_0671_),
    .A2(_0675_),
    .B(\Control_unit1.instr_stage1[0] ),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2830_ (.A1(_0616_),
    .A2(_2086_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2831_ (.I(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2832_ (.A1(_2079_),
    .A2(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2833_ (.A1(_0633_),
    .A2(_0676_),
    .A3(_0679_),
    .ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2834_ (.I(_0677_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2835_ (.A1(_2084_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2836_ (.I(_0670_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2837_ (.I(_0618_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2838_ (.A1(_0616_),
    .A2(_0683_),
    .B(_0674_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2839_ (.I(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2840_ (.A1(\Control_unit1.instr_stage1[1] ),
    .A2(_0682_),
    .B1(_0685_),
    .B2(\Stack_pointer.SP[1] ),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2841_ (.A1(_0681_),
    .A2(_0686_),
    .ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2842_ (.I(_2101_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2843_ (.I(_0687_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2844_ (.A1(_0688_),
    .A2(_0678_),
    .B1(_0671_),
    .B2(\Control_unit1.instr_stage1[2] ),
    .C1(_0684_),
    .C2(\Stack_pointer.SP[2] ),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2845_ (.I(_0689_),
    .ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2846_ (.A1(\Control_unit2.instr_stage2[3] ),
    .A2(_0680_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2847_ (.A1(\Control_unit1.instr_stage1[3] ),
    .A2(_0682_),
    .B1(_0685_),
    .B2(\Stack_pointer.SP[3] ),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2848_ (.A1(_0690_),
    .A2(_0691_),
    .ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2849_ (.A1(\Control_unit2.instr_stage2[4] ),
    .A2(_0680_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2850_ (.A1(\Control_unit1.instr_stage1[4] ),
    .A2(_0682_),
    .B1(_0685_),
    .B2(\Stack_pointer.SP[4] ),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2851_ (.A1(_0692_),
    .A2(_0693_),
    .ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2852_ (.A1(\Control_unit2.instr_stage2[5] ),
    .A2(_0680_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2853_ (.A1(\Control_unit1.instr_stage1[5] ),
    .A2(_0682_),
    .B1(_0685_),
    .B2(\Stack_pointer.SP[5] ),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2854_ (.A1(_0694_),
    .A2(_0695_),
    .ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2855_ (.A1(\Control_unit2.instr_stage2[6] ),
    .A2(_0678_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2856_ (.A1(\Control_unit1.instr_stage1[6] ),
    .A2(_0671_),
    .B1(_0684_),
    .B2(\Stack_pointer.SP[6] ),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2857_ (.A1(_0696_),
    .A2(_0697_),
    .ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2858_ (.A1(\Control_unit2.instr_stage2[7] ),
    .A2(_0678_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2859_ (.A1(\Control_unit1.instr_stage1[7] ),
    .A2(_0671_),
    .B1(_0684_),
    .B2(\Stack_pointer.SP[7] ),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2860_ (.A1(_0698_),
    .A2(_0699_),
    .ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2861_ (.I(\Control_unit2.instr_stage2[12] ),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2862_ (.I(\Arithmetic_Logic_Unit.ALU_001.p_Z ),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2863_ (.A1(_0700_),
    .A2(\Control_unit2.instr_stage2[11] ),
    .B(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2864_ (.I(\Control_unit2.instr_stage2[11] ),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2865_ (.A1(_2089_),
    .A2(_0703_),
    .B(\Arithmetic_Logic_Unit.ALU_001.p_Z ),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2866_ (.A1(_2088_),
    .A2(_0702_),
    .A3(_0704_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2867_ (.I(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2868_ (.A1(net70),
    .A2(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2869_ (.A1(_2088_),
    .A2(_2090_),
    .B(net35),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2870_ (.I(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2871_ (.I(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2872_ (.I(_0683_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2873_ (.I(_0711_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2874_ (.A1(_0683_),
    .A2(_0705_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2875_ (.I(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2876_ (.A1(net47),
    .A2(net51),
    .A3(net52),
    .A4(net53),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2877_ (.A1(net54),
    .A2(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2878_ (.A1(\Control_unit2.instr_stage2[4] ),
    .A2(_0712_),
    .B1(_0714_),
    .B2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2879_ (.A1(net35),
    .A2(net46),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2880_ (.I(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2881_ (.I(net54),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2882_ (.A1(_0707_),
    .A2(_0710_),
    .A3(_0717_),
    .B1(_0719_),
    .B2(_0720_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2883_ (.I(_0709_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2884_ (.A1(net54),
    .A2(_0715_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2885_ (.A1(net55),
    .A2(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2886_ (.A1(net55),
    .A2(_0722_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2887_ (.A1(_0723_),
    .A2(_0724_),
    .B(_0714_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2888_ (.I(_0705_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2889_ (.A1(\Control_unit2.instr_stage2[5] ),
    .A2(_0712_),
    .B1(_0726_),
    .B2(_2274_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2890_ (.I(net55),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2891_ (.A1(_0721_),
    .A2(_0725_),
    .A3(_0727_),
    .B1(_0719_),
    .B2(_0728_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2892_ (.I(net56),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2893_ (.I(_0718_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2894_ (.A1(_0683_),
    .A2(_0705_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2895_ (.I(_0731_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2896_ (.A1(net56),
    .A2(_0723_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2897_ (.A1(_0732_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2898_ (.A1(\Control_unit2.instr_stage2[6] ),
    .A2(_0712_),
    .B1(_0706_),
    .B2(_2250_),
    .C(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2899_ (.A1(_0729_),
    .A2(_0730_),
    .B1(_0710_),
    .B2(_0735_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2900_ (.I(net57),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2901_ (.A1(net55),
    .A2(net56),
    .A3(_0722_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2902_ (.A1(net57),
    .A2(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2903_ (.A1(_0731_),
    .A2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2904_ (.A1(\Control_unit2.instr_stage2[7] ),
    .A2(_0712_),
    .B1(_0706_),
    .B2(_2273_),
    .C(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2905_ (.A1(_0736_),
    .A2(_0719_),
    .B1(_0710_),
    .B2(_0740_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2906_ (.A1(_0736_),
    .A2(_0737_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2907_ (.A1(net58),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2908_ (.I(net58),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2909_ (.A1(_0736_),
    .A2(_0737_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2910_ (.A1(_0742_),
    .A2(_0744_),
    .B(_0714_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2911_ (.I(\Control_unit2.instr_stage2[8] ),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2912_ (.I(_0711_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2913_ (.A1(_0746_),
    .A2(_0747_),
    .B1(_0726_),
    .B2(_2283_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2914_ (.I(_0718_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2915_ (.A1(_0721_),
    .A2(_0745_),
    .A3(_0748_),
    .B1(_0749_),
    .B2(_0743_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2916_ (.I(net59),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2917_ (.I(\Control_unit2.instr_stage2[9] ),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2918_ (.A1(_2088_),
    .A2(_0702_),
    .A3(_0704_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2919_ (.I(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2920_ (.A1(net59),
    .A2(_0742_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2921_ (.A1(_2335_),
    .A2(_0753_),
    .B1(_0732_),
    .B2(_0754_),
    .C(_0709_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2922_ (.A1(_0751_),
    .A2(_0667_),
    .B(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2923_ (.A1(_0750_),
    .A2(_0730_),
    .B(_0756_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2924_ (.A1(_2341_),
    .A2(_2353_),
    .B(_0726_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2925_ (.I(\Control_unit2.instr_stage2[10] ),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2926_ (.I(net48),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2927_ (.A1(net58),
    .A2(net59),
    .A3(_0741_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2928_ (.A1(_0759_),
    .A2(_0760_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2929_ (.A1(_0758_),
    .A2(_0747_),
    .B1(_0714_),
    .B2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2930_ (.A1(_0721_),
    .A2(_0757_),
    .A3(_0762_),
    .B1(_0749_),
    .B2(_0759_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2931_ (.A1(net62),
    .A2(_0706_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2932_ (.I(\Control_unit2.instr_stage2[11] ),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2933_ (.A1(_0759_),
    .A2(_0760_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2934_ (.A1(net49),
    .A2(_0765_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2935_ (.A1(_0764_),
    .A2(_0747_),
    .B1(_0713_),
    .B2(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2936_ (.I(net49),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2937_ (.A1(_0721_),
    .A2(_0763_),
    .A3(_0767_),
    .B1(_0749_),
    .B2(_0768_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2938_ (.I(net50),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2939_ (.A1(net49),
    .A2(_0765_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2940_ (.A1(net50),
    .A2(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2941_ (.A1(_0711_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2942_ (.A1(_2089_),
    .A2(_0711_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2943_ (.I0(_0571_),
    .I1(_0773_),
    .S(_0726_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2944_ (.A1(_0769_),
    .A2(_0719_),
    .B1(_0710_),
    .B2(_0774_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2945_ (.A1(\Control_unit1.instr_stage1[0] ),
    .A2(_0673_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2946_ (.A1(_0624_),
    .A2(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2947_ (.A1(_0669_),
    .A2(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2948_ (.I(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2949_ (.I(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2950_ (.I(net18),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2951_ (.I(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2952_ (.I(_0777_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2953_ (.I(_0782_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2954_ (.A1(_0781_),
    .A2(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2955_ (.A1(_2146_),
    .A2(_0779_),
    .B(_0784_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2956_ (.I(net25),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2957_ (.I(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2958_ (.A1(_0786_),
    .A2(_0783_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2959_ (.A1(_2172_),
    .A2(_0779_),
    .B(_0787_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2960_ (.I(net26),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2961_ (.I(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2962_ (.A1(_0789_),
    .A2(_0783_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2963_ (.A1(_2190_),
    .A2(_0779_),
    .B(_0790_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2964_ (.I(net27),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2965_ (.I(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2966_ (.A1(_0792_),
    .A2(_0783_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2967_ (.A1(_2212_),
    .A2(_0779_),
    .B(_0793_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2968_ (.I(_2232_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2969_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2970_ (.I(_0778_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2971_ (.I(net28),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2972_ (.I(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2973_ (.I(_0782_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2974_ (.A1(_0798_),
    .A2(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2975_ (.A1(_0795_),
    .A2(_0796_),
    .B(_0800_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2976_ (.I(net29),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2977_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2978_ (.A1(_0802_),
    .A2(_0799_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2979_ (.A1(_2257_),
    .A2(_0796_),
    .B(_0803_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2980_ (.I(net30),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2981_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2982_ (.A1(_0805_),
    .A2(_0799_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2983_ (.A1(_2278_),
    .A2(_0796_),
    .B(_0806_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2984_ (.I(net31),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2985_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2986_ (.A1(_0808_),
    .A2(_0799_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2987_ (.A1(_2298_),
    .A2(_0796_),
    .B(_0809_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2988_ (.I(_0778_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2989_ (.I(net32),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2990_ (.I(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2991_ (.I(_0782_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2992_ (.A1(_0812_),
    .A2(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2993_ (.A1(_2322_),
    .A2(_0810_),
    .B(_0814_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2994_ (.I(net33),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2995_ (.I(_0815_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2996_ (.A1(_0816_),
    .A2(_0813_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2997_ (.A1(_2336_),
    .A2(_0810_),
    .B(_0817_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2998_ (.I(net19),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2999_ (.I(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3000_ (.A1(_0819_),
    .A2(_0813_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3001_ (.A1(_2355_),
    .A2(_0810_),
    .B(_0820_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3002_ (.I(_2370_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3003_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3004_ (.I(net20),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3005_ (.I(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3006_ (.A1(_0824_),
    .A2(_0813_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3007_ (.A1(_0822_),
    .A2(_0810_),
    .B(_0825_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3008_ (.I(_0778_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3009_ (.I(net21),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3010_ (.I(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3011_ (.I(_0782_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3012_ (.A1(_0828_),
    .A2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3013_ (.A1(_0572_),
    .A2(_0826_),
    .B(_0830_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3014_ (.I(net22),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3015_ (.I(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3016_ (.A1(_0832_),
    .A2(_0829_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3017_ (.A1(_0592_),
    .A2(_0826_),
    .B(_0833_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3018_ (.I(net23),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3019_ (.I(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3020_ (.A1(_0835_),
    .A2(_0829_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3021_ (.A1(_0604_),
    .A2(_0826_),
    .B(_0836_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3022_ (.I(net24),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3023_ (.I(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3024_ (.A1(_0838_),
    .A2(_0829_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3025_ (.A1(_0615_),
    .A2(_0826_),
    .B(_0839_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3026_ (.A1(\Control_unit1.instr_decoder1.A[2] ),
    .A2(\Control_unit1.instr_decoder1.A[1] ),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3027_ (.A1(_0840_),
    .A2(_0623_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3028_ (.I(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3029_ (.I(_0842_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3030_ (.I(_0841_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3031_ (.A1(_0780_),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3032_ (.A1(_2097_),
    .A2(_0843_),
    .B(_0845_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3033_ (.A1(_0785_),
    .A2(_0844_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3034_ (.A1(_2151_),
    .A2(_0843_),
    .B(_0846_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3035_ (.A1(_0788_),
    .A2(_0844_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3036_ (.A1(_2177_),
    .A2(_0843_),
    .B(_0847_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3037_ (.I(_0841_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3038_ (.A1(_0791_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3039_ (.A1(_2193_),
    .A2(_0843_),
    .B(_0849_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3040_ (.I0(_0798_),
    .I1(_2206_),
    .S(_0848_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3041_ (.I(_0850_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3042_ (.I0(_0802_),
    .I1(_2274_),
    .S(_0848_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3043_ (.I(_0851_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3044_ (.I(_0842_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3045_ (.I0(_0805_),
    .I1(_2250_),
    .S(_0852_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3046_ (.I(_0853_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3047_ (.I0(_0808_),
    .I1(_2273_),
    .S(_0852_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3048_ (.I(_0854_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3049_ (.I0(_0812_),
    .I1(_2283_),
    .S(_0852_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3050_ (.I(_0855_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3051_ (.I0(_0816_),
    .I1(_2318_),
    .S(_0852_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3052_ (.I(_0856_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3053_ (.A1(_0818_),
    .A2(_0848_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3054_ (.A1(_2338_),
    .A2(_0844_),
    .B(_0857_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3055_ (.I(_0842_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3056_ (.I0(_0824_),
    .I1(_2337_),
    .S(_0858_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3057_ (.I(_0859_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3058_ (.I0(_0828_),
    .I1(_2366_),
    .S(_0858_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3059_ (.I(_0860_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3060_ (.I0(_0832_),
    .I1(_0567_),
    .S(_0858_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3061_ (.I(_0861_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3062_ (.I0(_0835_),
    .I1(_0588_),
    .S(_0858_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3063_ (.I(_0862_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3064_ (.I0(_0838_),
    .I1(_0612_),
    .S(_0842_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3065_ (.I(_0863_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3066_ (.A1(_0687_),
    .A2(_2233_),
    .B(\Control_unit2.instr_decoder2.A[2] ),
    .C(\Control_unit2.instr_decoder2.A[1] ),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3067_ (.I(_2233_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3068_ (.A1(_2106_),
    .A2(_2251_),
    .B1(_2253_),
    .B2(_0612_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3069_ (.A1(_0865_),
    .A2(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3070_ (.A1(_0864_),
    .A2(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3071_ (.I(_0610_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3072_ (.A1(_0608_),
    .A2(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3073_ (.A1(_0596_),
    .A2(_0606_),
    .B(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3074_ (.A1(_0584_),
    .A2(_0605_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3075_ (.A1(_0612_),
    .A2(_2261_),
    .A3(_0610_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3076_ (.A1(_0872_),
    .A2(_0873_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3077_ (.A1(_0871_),
    .A2(_0874_),
    .B(_0688_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3078_ (.A1(_0688_),
    .A2(_0871_),
    .A3(_0874_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3079_ (.A1(_0865_),
    .A2(_0875_),
    .A3(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3080_ (.A1(_2121_),
    .A2(_0864_),
    .B1(_0868_),
    .B2(_0877_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3081_ (.A1(\Control_unit2.instr_stage2[9] ),
    .A2(\Control_unit2.instr_stage2[10] ),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3082_ (.A1(_0746_),
    .A2(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3083_ (.A1(_0687_),
    .A2(\Control_unit2.instr_decoder2.A[1] ),
    .B(_2141_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3084_ (.A1(_2119_),
    .A2(_2087_),
    .B1(_0880_),
    .B2(_2085_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3085_ (.A1(_0700_),
    .A2(_0764_),
    .A3(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3086_ (.I(_0882_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3087_ (.A1(_0879_),
    .A2(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3088_ (.I(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3089_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3090_ (.I(_0884_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3091_ (.I(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3092_ (.A1(_0781_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3093_ (.A1(_2146_),
    .A2(_0886_),
    .B(_0889_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3094_ (.A1(_0786_),
    .A2(_0888_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3095_ (.A1(_2172_),
    .A2(_0886_),
    .B(_0890_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3096_ (.A1(_0789_),
    .A2(_0888_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3097_ (.A1(_2190_),
    .A2(_0886_),
    .B(_0891_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3098_ (.A1(_0792_),
    .A2(_0888_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3099_ (.A1(_2212_),
    .A2(_0886_),
    .B(_0892_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3100_ (.I(_0885_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3101_ (.I(_0887_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3102_ (.A1(_0798_),
    .A2(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3103_ (.A1(_0795_),
    .A2(_0893_),
    .B(_0895_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3104_ (.A1(_0802_),
    .A2(_0894_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3105_ (.A1(_2257_),
    .A2(_0893_),
    .B(_0896_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3106_ (.A1(_0805_),
    .A2(_0894_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3107_ (.A1(_2278_),
    .A2(_0893_),
    .B(_0897_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3108_ (.A1(_0808_),
    .A2(_0894_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3109_ (.A1(_2298_),
    .A2(_0893_),
    .B(_0898_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3110_ (.I(_0885_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3111_ (.I(_0887_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3112_ (.A1(_0812_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3113_ (.A1(_2322_),
    .A2(_0899_),
    .B(_0901_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3114_ (.A1(_0816_),
    .A2(_0900_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3115_ (.A1(_2336_),
    .A2(_0899_),
    .B(_0902_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3116_ (.A1(_0819_),
    .A2(_0900_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3117_ (.A1(_2355_),
    .A2(_0899_),
    .B(_0903_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3118_ (.A1(_0824_),
    .A2(_0900_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3119_ (.A1(_0822_),
    .A2(_0899_),
    .B(_0904_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3120_ (.I(_0885_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3121_ (.I(_0887_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3122_ (.A1(_0828_),
    .A2(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3123_ (.A1(_0572_),
    .A2(_0905_),
    .B(_0907_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3124_ (.A1(_0832_),
    .A2(_0906_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3125_ (.A1(_0592_),
    .A2(_0905_),
    .B(_0908_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3126_ (.A1(_0835_),
    .A2(_0906_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3127_ (.A1(_0604_),
    .A2(_0905_),
    .B(_0909_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3128_ (.A1(_0838_),
    .A2(_0906_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3129_ (.A1(_0615_),
    .A2(_0905_),
    .B(_0910_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3130_ (.A1(_2349_),
    .A2(_2352_),
    .B1(_0561_),
    .B2(_0564_),
    .C(_2332_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3131_ (.A1(_2312_),
    .A2(_2313_),
    .B(_2314_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3132_ (.A1(_2300_),
    .A2(_2303_),
    .A3(_2309_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3133_ (.A1(_2241_),
    .A2(_2246_),
    .B1(_2269_),
    .B2(_2270_),
    .C1(_0912_),
    .C2(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3134_ (.A1(_0687_),
    .A2(_2251_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3135_ (.A1(_2129_),
    .A2(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3136_ (.A1(_2161_),
    .A2(_2183_),
    .A3(_2228_),
    .A4(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3137_ (.A1(_2204_),
    .A2(_2295_),
    .A3(_0914_),
    .A4(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3138_ (.A1(_2364_),
    .A2(_0585_),
    .A3(_0911_),
    .A4(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3139_ (.A1(_0600_),
    .A2(_0919_),
    .B(_0865_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3140_ (.A1(_2206_),
    .A2(_2274_),
    .A3(_2250_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3141_ (.A1(_2084_),
    .A2(_2135_),
    .A3(_2165_),
    .A4(_2185_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3142_ (.A1(_0921_),
    .A2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3143_ (.A1(_2319_),
    .A2(_2333_),
    .A3(_2340_),
    .A4(_2368_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3144_ (.A1(_2285_),
    .A2(_0923_),
    .A3(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3145_ (.A1(_0568_),
    .A2(_0589_),
    .A3(_0602_),
    .A4(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3146_ (.A1(_2140_),
    .A2(_0613_),
    .A3(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3147_ (.A1(_0586_),
    .A2(_0701_),
    .B(_0927_),
    .C(_2233_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3148_ (.A1(_0865_),
    .A2(_0611_),
    .B(_0864_),
    .C(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3149_ (.A1(_0701_),
    .A2(_0864_),
    .B1(_0920_),
    .B2(_0929_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3150_ (.I(\Control_unit2.instr_stage2[8] ),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3151_ (.A1(_0930_),
    .A2(\Control_unit2.instr_stage2[9] ),
    .A3(\Control_unit2.instr_stage2[10] ),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3152_ (.A1(_2089_),
    .A2(_0764_),
    .A3(_0881_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3153_ (.I(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3154_ (.A1(_0931_),
    .A2(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3155_ (.I(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3156_ (.I(_0935_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3157_ (.I(_0934_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3158_ (.I(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3159_ (.A1(_0781_),
    .A2(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3160_ (.A1(_2146_),
    .A2(_0936_),
    .B(_0939_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3161_ (.A1(_0786_),
    .A2(_0938_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3162_ (.A1(_2172_),
    .A2(_0936_),
    .B(_0940_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3163_ (.A1(_0789_),
    .A2(_0938_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3164_ (.A1(_2190_),
    .A2(_0936_),
    .B(_0941_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3165_ (.A1(_0792_),
    .A2(_0938_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3166_ (.A1(_2212_),
    .A2(_0936_),
    .B(_0942_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3167_ (.I(_0935_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3168_ (.I(_0937_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3169_ (.A1(_0798_),
    .A2(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3170_ (.A1(_0795_),
    .A2(_0943_),
    .B(_0945_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3171_ (.A1(_0802_),
    .A2(_0944_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3172_ (.A1(_2257_),
    .A2(_0943_),
    .B(_0946_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3173_ (.A1(_0805_),
    .A2(_0944_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3174_ (.A1(_2278_),
    .A2(_0943_),
    .B(_0947_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3175_ (.A1(_0808_),
    .A2(_0944_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3176_ (.A1(_2298_),
    .A2(_0943_),
    .B(_0948_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3177_ (.I(_0935_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3178_ (.I(_0937_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3179_ (.A1(_0812_),
    .A2(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3180_ (.A1(_2322_),
    .A2(_0949_),
    .B(_0951_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3181_ (.A1(_0816_),
    .A2(_0950_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3182_ (.A1(_2336_),
    .A2(_0949_),
    .B(_0952_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3183_ (.A1(_0819_),
    .A2(_0950_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3184_ (.A1(_2355_),
    .A2(_0949_),
    .B(_0953_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3185_ (.A1(_0824_),
    .A2(_0950_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3186_ (.A1(_0822_),
    .A2(_0949_),
    .B(_0954_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3187_ (.I(_0935_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3188_ (.I(_0937_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3189_ (.A1(_0828_),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3190_ (.A1(_0572_),
    .A2(_0955_),
    .B(_0957_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3191_ (.A1(_0832_),
    .A2(_0956_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3192_ (.A1(_0592_),
    .A2(_0955_),
    .B(_0958_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3193_ (.A1(_0835_),
    .A2(_0956_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3194_ (.A1(_0604_),
    .A2(_0955_),
    .B(_0959_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3195_ (.A1(_0838_),
    .A2(_0956_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3196_ (.A1(_0615_),
    .A2(_0955_),
    .B(_0960_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3197_ (.I(_2145_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3198_ (.I(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3199_ (.I(\Control_unit2.instr_stage2[10] ),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3200_ (.A1(_0930_),
    .A2(_0751_),
    .A3(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3201_ (.A1(_2090_),
    .A2(_0881_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3202_ (.I(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3203_ (.A1(_0964_),
    .A2(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3204_ (.I(_0967_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3205_ (.I(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3206_ (.I(_0967_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3207_ (.I(_0970_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3208_ (.A1(_0781_),
    .A2(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3209_ (.A1(_0962_),
    .A2(_0969_),
    .B(_0972_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3210_ (.I(_2171_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3211_ (.I(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3212_ (.A1(_0786_),
    .A2(_0971_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3213_ (.A1(_0974_),
    .A2(_0969_),
    .B(_0975_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3214_ (.I(_2189_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3215_ (.I(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3216_ (.A1(_0789_),
    .A2(_0971_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3217_ (.A1(_0977_),
    .A2(_0969_),
    .B(_0978_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3218_ (.I(_2211_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3219_ (.I(_0979_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3220_ (.A1(_0792_),
    .A2(_0971_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3221_ (.A1(_0980_),
    .A2(_0969_),
    .B(_0981_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3222_ (.I(_0968_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3223_ (.I(_0797_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3224_ (.I(_0970_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3225_ (.A1(_0983_),
    .A2(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3226_ (.A1(_0795_),
    .A2(_0982_),
    .B(_0985_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3227_ (.I(_2256_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3228_ (.I(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3229_ (.I(_0801_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3230_ (.A1(_0988_),
    .A2(_0984_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3231_ (.A1(_0987_),
    .A2(_0982_),
    .B(_0989_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3232_ (.I(_2277_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3233_ (.I(_0990_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3234_ (.I(_0804_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3235_ (.A1(_0992_),
    .A2(_0984_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3236_ (.A1(_0991_),
    .A2(_0982_),
    .B(_0993_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3237_ (.I(_2297_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3238_ (.I(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3239_ (.I(_0807_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3240_ (.A1(_0996_),
    .A2(_0984_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3241_ (.A1(_0995_),
    .A2(_0982_),
    .B(_0997_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3242_ (.I(_2321_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3243_ (.I(_0998_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3244_ (.I(_0968_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3245_ (.I(_0811_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3246_ (.I(_0970_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3247_ (.A1(_1001_),
    .A2(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3248_ (.A1(_0999_),
    .A2(_1000_),
    .B(_1003_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3249_ (.I(_2335_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3250_ (.I(_1004_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3251_ (.I(_0815_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3252_ (.A1(_1006_),
    .A2(_1002_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3253_ (.A1(_1005_),
    .A2(_1000_),
    .B(_1007_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3254_ (.I(_2354_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3255_ (.I(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3256_ (.A1(_0819_),
    .A2(_1002_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3257_ (.A1(_1009_),
    .A2(_1000_),
    .B(_1010_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3258_ (.I(_0823_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3259_ (.A1(_1011_),
    .A2(_1002_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3260_ (.A1(_0822_),
    .A2(_1000_),
    .B(_1012_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3261_ (.I(_0571_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3262_ (.I(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3263_ (.I(_0968_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3264_ (.I(_0827_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3265_ (.I(_0970_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3266_ (.A1(_1016_),
    .A2(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3267_ (.A1(_1014_),
    .A2(_1015_),
    .B(_1018_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3268_ (.I(_0591_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3269_ (.I(_1019_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3270_ (.I(_0831_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3271_ (.A1(_1021_),
    .A2(_1017_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3272_ (.A1(_1020_),
    .A2(_1015_),
    .B(_1022_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3273_ (.I(_0603_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3274_ (.I(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3275_ (.I(_0834_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3276_ (.A1(_1025_),
    .A2(_1017_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3277_ (.A1(_1024_),
    .A2(_1015_),
    .B(_1026_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3278_ (.I(_0614_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3279_ (.I(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3280_ (.I(_0837_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3281_ (.A1(_1029_),
    .A2(_1017_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3282_ (.A1(_1028_),
    .A2(_1015_),
    .B(_1030_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3283_ (.I(_0932_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3284_ (.I(\Control_unit2.instr_stage2[9] ),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3285_ (.A1(_0930_),
    .A2(_1032_),
    .A3(_0758_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3286_ (.A1(_1031_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3287_ (.I(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3288_ (.I(_1035_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3289_ (.I(_0780_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3290_ (.I(_1034_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3291_ (.I(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3292_ (.A1(_1037_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3293_ (.A1(_0962_),
    .A2(_1036_),
    .B(_1040_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3294_ (.I(_0785_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3295_ (.A1(_1041_),
    .A2(_1039_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3296_ (.A1(_0974_),
    .A2(_1036_),
    .B(_1042_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3297_ (.I(_0788_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3298_ (.A1(_1043_),
    .A2(_1039_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3299_ (.A1(_0977_),
    .A2(_1036_),
    .B(_1044_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3300_ (.I(_0791_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3301_ (.A1(_1045_),
    .A2(_1039_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3302_ (.A1(_0980_),
    .A2(_1036_),
    .B(_1046_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3303_ (.I(_0794_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3304_ (.I(_1035_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3305_ (.I(_1038_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3306_ (.A1(_0983_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3307_ (.A1(_1047_),
    .A2(_1048_),
    .B(_1050_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3308_ (.A1(_0988_),
    .A2(_1049_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3309_ (.A1(_0987_),
    .A2(_1048_),
    .B(_1051_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3310_ (.A1(_0992_),
    .A2(_1049_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3311_ (.A1(_0991_),
    .A2(_1048_),
    .B(_1052_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3312_ (.A1(_0996_),
    .A2(_1049_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3313_ (.A1(_0995_),
    .A2(_1048_),
    .B(_1053_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3314_ (.I(_1035_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3315_ (.I(_1038_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3316_ (.A1(_1001_),
    .A2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3317_ (.A1(_0999_),
    .A2(_1054_),
    .B(_1056_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3318_ (.A1(_1006_),
    .A2(_1055_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3319_ (.A1(_1005_),
    .A2(_1054_),
    .B(_1057_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3320_ (.I(_0818_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3321_ (.A1(_1058_),
    .A2(_1055_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3322_ (.A1(_1009_),
    .A2(_1054_),
    .B(_1059_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3323_ (.I(_0821_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3324_ (.A1(_1011_),
    .A2(_1055_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3325_ (.A1(_1060_),
    .A2(_1054_),
    .B(_1061_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3326_ (.I(_1035_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3327_ (.I(_1038_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3328_ (.A1(_1016_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3329_ (.A1(_1014_),
    .A2(_1062_),
    .B(_1064_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3330_ (.A1(_1021_),
    .A2(_1063_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3331_ (.A1(_1020_),
    .A2(_1062_),
    .B(_1065_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3332_ (.A1(_1025_),
    .A2(_1063_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3333_ (.A1(_1024_),
    .A2(_1062_),
    .B(_1066_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3334_ (.A1(_1029_),
    .A2(_1063_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3335_ (.A1(_1028_),
    .A2(_1062_),
    .B(_1067_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3336_ (.A1(_0746_),
    .A2(_0751_),
    .A3(_0963_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3337_ (.A1(_1031_),
    .A2(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3338_ (.I(_1069_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3339_ (.I(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3340_ (.I(_1069_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3341_ (.I(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3342_ (.A1(_1037_),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3343_ (.A1(_0962_),
    .A2(_1071_),
    .B(_1074_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3344_ (.A1(_1041_),
    .A2(_1073_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3345_ (.A1(_0974_),
    .A2(_1071_),
    .B(_1075_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3346_ (.A1(_1043_),
    .A2(_1073_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3347_ (.A1(_0977_),
    .A2(_1071_),
    .B(_1076_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3348_ (.A1(_1045_),
    .A2(_1073_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3349_ (.A1(_0980_),
    .A2(_1071_),
    .B(_1077_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3350_ (.I(_1070_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3351_ (.I(_1072_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3352_ (.A1(_0983_),
    .A2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3353_ (.A1(_1047_),
    .A2(_1078_),
    .B(_1080_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3354_ (.A1(_0988_),
    .A2(_1079_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3355_ (.A1(_0987_),
    .A2(_1078_),
    .B(_1081_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3356_ (.A1(_0992_),
    .A2(_1079_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3357_ (.A1(_0991_),
    .A2(_1078_),
    .B(_1082_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3358_ (.A1(_0996_),
    .A2(_1079_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3359_ (.A1(_0995_),
    .A2(_1078_),
    .B(_1083_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3360_ (.I(_1070_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3361_ (.I(_1072_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3362_ (.A1(_1001_),
    .A2(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3363_ (.A1(_0999_),
    .A2(_1084_),
    .B(_1086_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3364_ (.A1(_1006_),
    .A2(_1085_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3365_ (.A1(_1005_),
    .A2(_1084_),
    .B(_1087_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3366_ (.A1(_1058_),
    .A2(_1085_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3367_ (.A1(_1009_),
    .A2(_1084_),
    .B(_1088_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3368_ (.A1(_1011_),
    .A2(_1085_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3369_ (.A1(_1060_),
    .A2(_1084_),
    .B(_1089_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3370_ (.I(_1070_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3371_ (.I(_1072_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3372_ (.A1(_1016_),
    .A2(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3373_ (.A1(_1014_),
    .A2(_1090_),
    .B(_1092_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3374_ (.A1(_1021_),
    .A2(_1091_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3375_ (.A1(_1020_),
    .A2(_1090_),
    .B(_1093_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3376_ (.A1(_1025_),
    .A2(_1091_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3377_ (.A1(_1024_),
    .A2(_1090_),
    .B(_1094_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3378_ (.A1(_1029_),
    .A2(_1091_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3379_ (.A1(_1028_),
    .A2(_1090_),
    .B(_1095_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3380_ (.A1(_1031_),
    .A2(_0964_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3381_ (.I(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3382_ (.I(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3383_ (.I(_1096_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3384_ (.I(_1099_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3385_ (.A1(_1037_),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3386_ (.A1(_0962_),
    .A2(_1098_),
    .B(_1101_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3387_ (.A1(_1041_),
    .A2(_1100_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3388_ (.A1(_0974_),
    .A2(_1098_),
    .B(_1102_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3389_ (.A1(_1043_),
    .A2(_1100_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3390_ (.A1(_0977_),
    .A2(_1098_),
    .B(_1103_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3391_ (.A1(_1045_),
    .A2(_1100_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3392_ (.A1(_0980_),
    .A2(_1098_),
    .B(_1104_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3393_ (.I(_1097_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3394_ (.I(_1099_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3395_ (.A1(_0983_),
    .A2(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3396_ (.A1(_1047_),
    .A2(_1105_),
    .B(_1107_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3397_ (.A1(_0988_),
    .A2(_1106_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3398_ (.A1(_0987_),
    .A2(_1105_),
    .B(_1108_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3399_ (.A1(_0992_),
    .A2(_1106_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3400_ (.A1(_0991_),
    .A2(_1105_),
    .B(_1109_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3401_ (.A1(_0996_),
    .A2(_1106_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3402_ (.A1(_0995_),
    .A2(_1105_),
    .B(_1110_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3403_ (.I(_1097_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3404_ (.I(_1099_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3405_ (.A1(_1001_),
    .A2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3406_ (.A1(_0999_),
    .A2(_1111_),
    .B(_1113_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3407_ (.A1(_1006_),
    .A2(_1112_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3408_ (.A1(_1005_),
    .A2(_1111_),
    .B(_1114_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3409_ (.A1(_1058_),
    .A2(_1112_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3410_ (.A1(_1009_),
    .A2(_1111_),
    .B(_1115_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3411_ (.A1(_1011_),
    .A2(_1112_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3412_ (.A1(_1060_),
    .A2(_1111_),
    .B(_1116_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3413_ (.I(_1097_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3414_ (.I(_1099_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3415_ (.A1(_1016_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3416_ (.A1(_1014_),
    .A2(_1117_),
    .B(_1119_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3417_ (.A1(_1021_),
    .A2(_1118_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3418_ (.A1(_1020_),
    .A2(_1117_),
    .B(_1120_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3419_ (.A1(_1025_),
    .A2(_1118_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3420_ (.A1(_1024_),
    .A2(_1117_),
    .B(_1121_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3421_ (.A1(_1029_),
    .A2(_1118_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3422_ (.A1(_1028_),
    .A2(_1117_),
    .B(_1122_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3423_ (.I(_0961_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3424_ (.A1(_0879_),
    .A2(_0933_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3425_ (.I(_1124_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3426_ (.I(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3427_ (.I(_1124_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3428_ (.I(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3429_ (.A1(_1037_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3430_ (.A1(_1123_),
    .A2(_1126_),
    .B(_1129_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3431_ (.I(_0973_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3432_ (.A1(_1041_),
    .A2(_1128_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3433_ (.A1(_1130_),
    .A2(_1126_),
    .B(_1131_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3434_ (.I(_0976_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3435_ (.A1(_1043_),
    .A2(_1128_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3436_ (.A1(_1132_),
    .A2(_1126_),
    .B(_1133_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3437_ (.I(_0979_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3438_ (.A1(_1045_),
    .A2(_1128_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3439_ (.A1(_1134_),
    .A2(_1126_),
    .B(_1135_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3440_ (.I(_1125_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3441_ (.I(net28),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3442_ (.I(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3443_ (.I(_1127_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3444_ (.A1(_1138_),
    .A2(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3445_ (.A1(_1047_),
    .A2(_1136_),
    .B(_1140_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3446_ (.I(_0986_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3447_ (.I(net29),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3448_ (.I(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3449_ (.A1(_1143_),
    .A2(_1139_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3450_ (.A1(_1141_),
    .A2(_1136_),
    .B(_1144_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3451_ (.I(_0990_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3452_ (.I(net30),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3453_ (.I(_1146_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3454_ (.A1(_1147_),
    .A2(_1139_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3455_ (.A1(_1145_),
    .A2(_1136_),
    .B(_1148_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3456_ (.I(_0994_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3457_ (.I(net31),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3458_ (.I(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3459_ (.A1(_1151_),
    .A2(_1139_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3460_ (.A1(_1149_),
    .A2(_1136_),
    .B(_1152_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3461_ (.I(_0998_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3462_ (.I(_1125_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3463_ (.I(net32),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3464_ (.I(_1155_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3465_ (.I(_1127_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3466_ (.A1(_1156_),
    .A2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3467_ (.A1(_1153_),
    .A2(_1154_),
    .B(_1158_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3468_ (.I(_1004_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3469_ (.I(net33),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3470_ (.I(_1160_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3471_ (.A1(_1161_),
    .A2(_1157_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3472_ (.A1(_1159_),
    .A2(_1154_),
    .B(_1162_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3473_ (.I(_1008_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3474_ (.A1(_1058_),
    .A2(_1157_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3475_ (.A1(_1163_),
    .A2(_1154_),
    .B(_1164_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3476_ (.I(net20),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3477_ (.I(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3478_ (.A1(_1166_),
    .A2(_1157_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3479_ (.A1(_1060_),
    .A2(_1154_),
    .B(_1167_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3480_ (.I(_1013_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3481_ (.I(_1125_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3482_ (.I(net21),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3483_ (.I(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3484_ (.I(_1127_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3485_ (.A1(_1171_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3486_ (.A1(_1168_),
    .A2(_1169_),
    .B(_1173_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3487_ (.I(_1019_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3488_ (.I(net22),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3489_ (.I(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3490_ (.A1(_1176_),
    .A2(_1172_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3491_ (.A1(_1174_),
    .A2(_1169_),
    .B(_1177_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3492_ (.I(_1023_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3493_ (.I(net23),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3494_ (.I(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3495_ (.A1(_1180_),
    .A2(_1172_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3496_ (.A1(_1178_),
    .A2(_1169_),
    .B(_1181_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3497_ (.I(_1027_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3498_ (.I(net24),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3499_ (.I(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3500_ (.A1(_1184_),
    .A2(_1172_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3501_ (.A1(_1182_),
    .A2(_1169_),
    .B(_1185_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3502_ (.A1(_0930_),
    .A2(_0878_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3503_ (.A1(_1031_),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3504_ (.I(_1187_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3505_ (.I(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3506_ (.I(net18),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3507_ (.I(_1190_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3508_ (.I(_1187_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3509_ (.I(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3510_ (.A1(_1191_),
    .A2(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3511_ (.A1(_1123_),
    .A2(_1189_),
    .B(_1194_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3512_ (.I(net25),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3513_ (.I(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3514_ (.A1(_1196_),
    .A2(_1193_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3515_ (.A1(_1130_),
    .A2(_1189_),
    .B(_1197_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3516_ (.I(net26),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3517_ (.I(_1198_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3518_ (.A1(_1199_),
    .A2(_1193_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3519_ (.A1(_1132_),
    .A2(_1189_),
    .B(_1200_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3520_ (.I(net27),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3521_ (.I(_1201_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3522_ (.A1(_1202_),
    .A2(_1193_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3523_ (.A1(_1134_),
    .A2(_1189_),
    .B(_1203_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3524_ (.I(_0794_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3525_ (.I(_1188_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3526_ (.I(_1192_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3527_ (.A1(_1138_),
    .A2(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3528_ (.A1(_1204_),
    .A2(_1205_),
    .B(_1207_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3529_ (.A1(_1143_),
    .A2(_1206_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3530_ (.A1(_1141_),
    .A2(_1205_),
    .B(_1208_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3531_ (.A1(_1147_),
    .A2(_1206_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3532_ (.A1(_1145_),
    .A2(_1205_),
    .B(_1209_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3533_ (.A1(_1151_),
    .A2(_1206_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3534_ (.A1(_1149_),
    .A2(_1205_),
    .B(_1210_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3535_ (.I(_1188_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3536_ (.I(_1192_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3537_ (.A1(_1156_),
    .A2(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3538_ (.A1(_1153_),
    .A2(_1211_),
    .B(_1213_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3539_ (.A1(_1161_),
    .A2(_1212_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3540_ (.A1(_1159_),
    .A2(_1211_),
    .B(_1214_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3541_ (.I(net19),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3542_ (.I(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3543_ (.A1(_1216_),
    .A2(_1212_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3544_ (.A1(_1163_),
    .A2(_1211_),
    .B(_1217_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3545_ (.I(_0821_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3546_ (.A1(_1166_),
    .A2(_1212_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3547_ (.A1(_1218_),
    .A2(_1211_),
    .B(_1219_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3548_ (.I(_1188_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3549_ (.I(_1192_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3550_ (.A1(_1171_),
    .A2(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3551_ (.A1(_1168_),
    .A2(_1220_),
    .B(_1222_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3552_ (.A1(_1176_),
    .A2(_1221_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3553_ (.A1(_1174_),
    .A2(_1220_),
    .B(_1223_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3554_ (.A1(_1180_),
    .A2(_1221_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3555_ (.A1(_1178_),
    .A2(_1220_),
    .B(_1224_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3556_ (.A1(_1184_),
    .A2(_1221_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3557_ (.A1(_1182_),
    .A2(_1220_),
    .B(_1225_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3558_ (.A1(\Control_unit2.instr_stage2[8] ),
    .A2(_0751_),
    .A3(_0758_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3559_ (.A1(_0700_),
    .A2(_0764_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3560_ (.A1(_1227_),
    .A2(_0881_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3561_ (.I(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3562_ (.A1(_1226_),
    .A2(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3563_ (.I(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3564_ (.I(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3565_ (.I(_1230_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3566_ (.I(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3567_ (.A1(_1191_),
    .A2(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3568_ (.A1(_1123_),
    .A2(_1232_),
    .B(_1235_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3569_ (.A1(_1196_),
    .A2(_1234_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3570_ (.A1(_1130_),
    .A2(_1232_),
    .B(_1236_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3571_ (.A1(_1199_),
    .A2(_1234_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3572_ (.A1(_1132_),
    .A2(_1232_),
    .B(_1237_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3573_ (.A1(_1202_),
    .A2(_1234_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3574_ (.A1(_1134_),
    .A2(_1232_),
    .B(_1238_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3575_ (.I(_1231_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3576_ (.I(_1233_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3577_ (.A1(_1138_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3578_ (.A1(_1204_),
    .A2(_1239_),
    .B(_1241_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3579_ (.A1(_1143_),
    .A2(_1240_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3580_ (.A1(_1141_),
    .A2(_1239_),
    .B(_1242_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3581_ (.A1(_1147_),
    .A2(_1240_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3582_ (.A1(_1145_),
    .A2(_1239_),
    .B(_1243_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3583_ (.A1(_1151_),
    .A2(_1240_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3584_ (.A1(_1149_),
    .A2(_1239_),
    .B(_1244_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3585_ (.I(_1231_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3586_ (.I(_1233_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3587_ (.A1(_1156_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3588_ (.A1(_1153_),
    .A2(_1245_),
    .B(_1247_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3589_ (.A1(_1161_),
    .A2(_1246_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3590_ (.A1(_1159_),
    .A2(_1245_),
    .B(_1248_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3591_ (.A1(_1216_),
    .A2(_1246_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3592_ (.A1(_1163_),
    .A2(_1245_),
    .B(_1249_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3593_ (.A1(_1166_),
    .A2(_1246_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3594_ (.A1(_1218_),
    .A2(_1245_),
    .B(_1250_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3595_ (.I(_1231_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3596_ (.I(_1233_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3597_ (.A1(_1171_),
    .A2(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3598_ (.A1(_1168_),
    .A2(_1251_),
    .B(_1253_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3599_ (.A1(_1176_),
    .A2(_1252_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3600_ (.A1(_1174_),
    .A2(_1251_),
    .B(_1254_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3601_ (.A1(_1180_),
    .A2(_1252_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3602_ (.A1(_1178_),
    .A2(_1251_),
    .B(_1255_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3603_ (.A1(_1184_),
    .A2(_1252_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3604_ (.A1(_1182_),
    .A2(_1251_),
    .B(_1256_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3605_ (.A1(_0931_),
    .A2(_1229_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3606_ (.I(_1257_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3607_ (.I(_1258_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3608_ (.I(_1257_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3609_ (.I(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3610_ (.A1(_1191_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3611_ (.A1(_1123_),
    .A2(_1259_),
    .B(_1262_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3612_ (.A1(_1196_),
    .A2(_1261_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3613_ (.A1(_1130_),
    .A2(_1259_),
    .B(_1263_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3614_ (.A1(_1199_),
    .A2(_1261_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3615_ (.A1(_1132_),
    .A2(_1259_),
    .B(_1264_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3616_ (.A1(_1202_),
    .A2(_1261_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3617_ (.A1(_1134_),
    .A2(_1259_),
    .B(_1265_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3618_ (.I(_1258_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3619_ (.I(_1260_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3620_ (.A1(_1138_),
    .A2(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3621_ (.A1(_1204_),
    .A2(_1266_),
    .B(_1268_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3622_ (.A1(_1143_),
    .A2(_1267_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3623_ (.A1(_1141_),
    .A2(_1266_),
    .B(_1269_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3624_ (.A1(_1147_),
    .A2(_1267_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3625_ (.A1(_1145_),
    .A2(_1266_),
    .B(_1270_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3626_ (.A1(_1151_),
    .A2(_1267_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3627_ (.A1(_1149_),
    .A2(_1266_),
    .B(_1271_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3628_ (.I(_1258_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3629_ (.I(_1260_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3630_ (.A1(_1156_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3631_ (.A1(_1153_),
    .A2(_1272_),
    .B(_1274_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3632_ (.A1(_1161_),
    .A2(_1273_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3633_ (.A1(_1159_),
    .A2(_1272_),
    .B(_1275_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3634_ (.A1(_1216_),
    .A2(_1273_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3635_ (.A1(_1163_),
    .A2(_1272_),
    .B(_1276_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3636_ (.A1(_1166_),
    .A2(_1273_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3637_ (.A1(_1218_),
    .A2(_1272_),
    .B(_1277_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3638_ (.I(_1258_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3639_ (.I(_1260_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3640_ (.A1(_1171_),
    .A2(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3641_ (.A1(_1168_),
    .A2(_1278_),
    .B(_1280_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3642_ (.A1(_1176_),
    .A2(_1279_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3643_ (.A1(_1174_),
    .A2(_1278_),
    .B(_1281_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3644_ (.A1(_1180_),
    .A2(_1279_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3645_ (.A1(_1178_),
    .A2(_1278_),
    .B(_1282_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3646_ (.A1(_1184_),
    .A2(_1279_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3647_ (.A1(_1182_),
    .A2(_1278_),
    .B(_1283_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3648_ (.I(_2144_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3649_ (.I(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3650_ (.A1(_0746_),
    .A2(_1032_),
    .A3(_0758_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3651_ (.A1(_1229_),
    .A2(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3652_ (.I(_1287_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3653_ (.I(_1288_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3654_ (.I(_1287_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3655_ (.I(_1290_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3656_ (.A1(_1191_),
    .A2(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3657_ (.A1(_1285_),
    .A2(_1289_),
    .B(_1292_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3658_ (.I(_2170_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3659_ (.I(_1293_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3660_ (.A1(_1196_),
    .A2(_1291_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3661_ (.A1(_1294_),
    .A2(_1289_),
    .B(_1295_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3662_ (.I(_2188_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3663_ (.I(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3664_ (.A1(_1199_),
    .A2(_1291_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3665_ (.A1(_1297_),
    .A2(_1289_),
    .B(_1298_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3666_ (.I(_2210_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3667_ (.I(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3668_ (.A1(_1202_),
    .A2(_1291_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3669_ (.A1(_1300_),
    .A2(_1289_),
    .B(_1301_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3670_ (.I(_1288_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3671_ (.I(_1137_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3672_ (.I(_1290_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3673_ (.A1(_1303_),
    .A2(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3674_ (.A1(_1204_),
    .A2(_1302_),
    .B(_1305_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3675_ (.I(_2256_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3676_ (.I(_1306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3677_ (.I(_1142_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3678_ (.A1(_1308_),
    .A2(_1304_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3679_ (.A1(_1307_),
    .A2(_1302_),
    .B(_1309_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3680_ (.I(_2277_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3681_ (.I(_1310_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3682_ (.I(_1146_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3683_ (.A1(_1312_),
    .A2(_1304_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3684_ (.A1(_1311_),
    .A2(_1302_),
    .B(_1313_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3685_ (.I(_2297_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3686_ (.I(_1314_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3687_ (.I(_1150_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3688_ (.A1(_1316_),
    .A2(_1304_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3689_ (.A1(_1315_),
    .A2(_1302_),
    .B(_1317_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3690_ (.I(_2321_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3691_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3692_ (.I(_1288_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3693_ (.I(_1155_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3694_ (.I(_1290_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3695_ (.A1(_1321_),
    .A2(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3696_ (.A1(_1319_),
    .A2(_1320_),
    .B(_1323_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3697_ (.I(_2334_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3698_ (.I(_1324_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3699_ (.I(_1160_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3700_ (.A1(_1326_),
    .A2(_1322_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3701_ (.A1(_1325_),
    .A2(_1320_),
    .B(_1327_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3702_ (.I(_2354_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3703_ (.I(_1328_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3704_ (.A1(_1216_),
    .A2(_1322_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3705_ (.A1(_1329_),
    .A2(_1320_),
    .B(_1330_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3706_ (.I(_1165_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3707_ (.A1(_1331_),
    .A2(_1322_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3708_ (.A1(_1218_),
    .A2(_1320_),
    .B(_1332_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3709_ (.I(_0570_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3710_ (.I(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3711_ (.I(_1288_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3712_ (.I(_1170_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3713_ (.I(_1290_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3714_ (.A1(_1336_),
    .A2(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3715_ (.A1(_1334_),
    .A2(_1335_),
    .B(_1338_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3716_ (.I(_0591_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3717_ (.I(_1339_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3718_ (.I(_1175_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3719_ (.A1(_1341_),
    .A2(_1337_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3720_ (.A1(_1340_),
    .A2(_1335_),
    .B(_1342_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3721_ (.I(_0603_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3722_ (.I(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3723_ (.I(_1179_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3724_ (.A1(_1345_),
    .A2(_1337_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3725_ (.A1(_1344_),
    .A2(_1335_),
    .B(_1346_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3726_ (.I(_0614_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3727_ (.I(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3728_ (.I(_1183_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3729_ (.A1(_1349_),
    .A2(_1337_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3730_ (.A1(_1348_),
    .A2(_1335_),
    .B(_1350_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3731_ (.A1(_1033_),
    .A2(_1229_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3732_ (.I(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3733_ (.I(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3734_ (.I(_1190_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3735_ (.I(_1351_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3736_ (.I(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3737_ (.A1(_1354_),
    .A2(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3738_ (.A1(_1285_),
    .A2(_1353_),
    .B(_1357_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3739_ (.I(_1195_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3740_ (.A1(_1358_),
    .A2(_1356_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3741_ (.A1(_1294_),
    .A2(_1353_),
    .B(_1359_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3742_ (.I(_1198_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3743_ (.A1(_1360_),
    .A2(_1356_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3744_ (.A1(_1297_),
    .A2(_1353_),
    .B(_1361_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3745_ (.I(_1201_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3746_ (.A1(_1362_),
    .A2(_1356_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3747_ (.A1(_1300_),
    .A2(_1353_),
    .B(_1363_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3748_ (.I(_2232_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3749_ (.I(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3750_ (.I(_1352_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3751_ (.I(_1355_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3752_ (.A1(_1303_),
    .A2(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3753_ (.A1(_1365_),
    .A2(_1366_),
    .B(_1368_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3754_ (.A1(_1308_),
    .A2(_1367_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3755_ (.A1(_1307_),
    .A2(_1366_),
    .B(_1369_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3756_ (.A1(_1312_),
    .A2(_1367_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3757_ (.A1(_1311_),
    .A2(_1366_),
    .B(_1370_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3758_ (.A1(_1316_),
    .A2(_1367_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3759_ (.A1(_1315_),
    .A2(_1366_),
    .B(_1371_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3760_ (.I(_1352_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3761_ (.I(_1355_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3762_ (.A1(_1321_),
    .A2(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3763_ (.A1(_1319_),
    .A2(_1372_),
    .B(_1374_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3764_ (.A1(_1326_),
    .A2(_1373_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3765_ (.A1(_1325_),
    .A2(_1372_),
    .B(_1375_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3766_ (.I(_1215_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3767_ (.A1(_1376_),
    .A2(_1373_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3768_ (.A1(_1329_),
    .A2(_1372_),
    .B(_1377_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3769_ (.I(_2370_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3770_ (.I(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3771_ (.A1(_1331_),
    .A2(_1373_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3772_ (.A1(_1379_),
    .A2(_1372_),
    .B(_1380_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3773_ (.I(_1352_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3774_ (.I(_1355_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3775_ (.A1(_1336_),
    .A2(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3776_ (.A1(_1334_),
    .A2(_1381_),
    .B(_1383_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3777_ (.A1(_1341_),
    .A2(_1382_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3778_ (.A1(_1340_),
    .A2(_1381_),
    .B(_1384_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3779_ (.A1(_1345_),
    .A2(_1382_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3780_ (.A1(_1344_),
    .A2(_1381_),
    .B(_1385_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3781_ (.A1(_1349_),
    .A2(_1382_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3782_ (.A1(_1348_),
    .A2(_1381_),
    .B(_1386_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3783_ (.A1(_0879_),
    .A2(_0966_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3784_ (.I(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3785_ (.I(_1388_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3786_ (.I(_1387_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3787_ (.I(_1390_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3788_ (.A1(_1354_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3789_ (.A1(_1285_),
    .A2(_1389_),
    .B(_1392_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3790_ (.A1(_1358_),
    .A2(_1391_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3791_ (.A1(_1294_),
    .A2(_1389_),
    .B(_1393_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3792_ (.A1(_1360_),
    .A2(_1391_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3793_ (.A1(_1297_),
    .A2(_1389_),
    .B(_1394_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3794_ (.A1(_1362_),
    .A2(_1391_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3795_ (.A1(_1300_),
    .A2(_1389_),
    .B(_1395_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3796_ (.I(_1388_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3797_ (.I(_1390_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3798_ (.A1(_1303_),
    .A2(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3799_ (.A1(_1365_),
    .A2(_1396_),
    .B(_1398_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3800_ (.A1(_1308_),
    .A2(_1397_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3801_ (.A1(_1307_),
    .A2(_1396_),
    .B(_1399_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3802_ (.A1(_1312_),
    .A2(_1397_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3803_ (.A1(_1311_),
    .A2(_1396_),
    .B(_1400_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3804_ (.A1(_1316_),
    .A2(_1397_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3805_ (.A1(_1315_),
    .A2(_1396_),
    .B(_1401_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3806_ (.I(_1388_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3807_ (.I(_1390_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3808_ (.A1(_1321_),
    .A2(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3809_ (.A1(_1319_),
    .A2(_1402_),
    .B(_1404_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3810_ (.A1(_1326_),
    .A2(_1403_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3811_ (.A1(_1325_),
    .A2(_1402_),
    .B(_1405_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3812_ (.A1(_1376_),
    .A2(_1403_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3813_ (.A1(_1329_),
    .A2(_1402_),
    .B(_1406_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3814_ (.A1(_1331_),
    .A2(_1403_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3815_ (.A1(_1379_),
    .A2(_1402_),
    .B(_1407_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3816_ (.I(_1388_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3817_ (.I(_1390_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3818_ (.A1(_1336_),
    .A2(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3819_ (.A1(_1334_),
    .A2(_1408_),
    .B(_1410_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3820_ (.A1(_1341_),
    .A2(_1409_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3821_ (.A1(_1340_),
    .A2(_1408_),
    .B(_1411_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3822_ (.A1(_1345_),
    .A2(_1409_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3823_ (.A1(_1344_),
    .A2(_1408_),
    .B(_1412_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3824_ (.A1(_1349_),
    .A2(_1409_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3825_ (.A1(_1348_),
    .A2(_1408_),
    .B(_1413_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3826_ (.I(_1228_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3827_ (.A1(_0964_),
    .A2(_1414_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3828_ (.I(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3829_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3830_ (.I(_1415_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3831_ (.I(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3832_ (.A1(_1354_),
    .A2(_1419_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3833_ (.A1(_1285_),
    .A2(_1417_),
    .B(_1420_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3834_ (.A1(_1358_),
    .A2(_1419_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3835_ (.A1(_1294_),
    .A2(_1417_),
    .B(_1421_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3836_ (.A1(_1360_),
    .A2(_1419_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3837_ (.A1(_1297_),
    .A2(_1417_),
    .B(_1422_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3838_ (.A1(_1362_),
    .A2(_1419_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3839_ (.A1(_1300_),
    .A2(_1417_),
    .B(_1423_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3840_ (.I(_1416_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3841_ (.I(_1418_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3842_ (.A1(_1303_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3843_ (.A1(_1365_),
    .A2(_1424_),
    .B(_1426_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3844_ (.A1(_1308_),
    .A2(_1425_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3845_ (.A1(_1307_),
    .A2(_1424_),
    .B(_1427_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3846_ (.A1(_1312_),
    .A2(_1425_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3847_ (.A1(_1311_),
    .A2(_1424_),
    .B(_1428_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3848_ (.A1(_1316_),
    .A2(_1425_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3849_ (.A1(_1315_),
    .A2(_1424_),
    .B(_1429_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3850_ (.I(_1416_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3851_ (.I(_1418_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3852_ (.A1(_1321_),
    .A2(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3853_ (.A1(_1319_),
    .A2(_1430_),
    .B(_1432_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3854_ (.A1(_1326_),
    .A2(_1431_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3855_ (.A1(_1325_),
    .A2(_1430_),
    .B(_1433_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3856_ (.A1(_1376_),
    .A2(_1431_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3857_ (.A1(_1329_),
    .A2(_1430_),
    .B(_1434_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3858_ (.A1(_1331_),
    .A2(_1431_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3859_ (.A1(_1379_),
    .A2(_1430_),
    .B(_1435_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3860_ (.I(_1416_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3861_ (.I(_1418_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3862_ (.A1(_1336_),
    .A2(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3863_ (.A1(_1334_),
    .A2(_1436_),
    .B(_1438_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3864_ (.A1(_1341_),
    .A2(_1437_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3865_ (.A1(_1340_),
    .A2(_1436_),
    .B(_1439_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3866_ (.A1(_1345_),
    .A2(_1437_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3867_ (.A1(_1344_),
    .A2(_1436_),
    .B(_1440_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3868_ (.A1(_1349_),
    .A2(_1437_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3869_ (.A1(_1348_),
    .A2(_1436_),
    .B(_1441_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3870_ (.I(_1284_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3871_ (.A1(_0879_),
    .A2(_1414_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3872_ (.I(_1443_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3873_ (.I(_1444_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3874_ (.I(_1443_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3875_ (.I(_1446_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3876_ (.A1(_1354_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3877_ (.A1(_1442_),
    .A2(_1445_),
    .B(_1448_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3878_ (.I(_1293_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3879_ (.A1(_1358_),
    .A2(_1447_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3880_ (.A1(_1449_),
    .A2(_1445_),
    .B(_1450_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3881_ (.I(_1296_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3882_ (.A1(_1360_),
    .A2(_1447_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3883_ (.A1(_1451_),
    .A2(_1445_),
    .B(_1452_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3884_ (.I(_1299_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3885_ (.A1(_1362_),
    .A2(_1447_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3886_ (.A1(_1453_),
    .A2(_1445_),
    .B(_1454_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3887_ (.I(_1444_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3888_ (.I(_1137_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3889_ (.I(_1446_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3890_ (.A1(_1456_),
    .A2(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3891_ (.A1(_1365_),
    .A2(_1455_),
    .B(_1458_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3892_ (.I(_1306_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3893_ (.I(_1142_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3894_ (.A1(_1460_),
    .A2(_1457_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3895_ (.A1(_1459_),
    .A2(_1455_),
    .B(_1461_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3896_ (.I(_1310_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3897_ (.I(_1146_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3898_ (.A1(_1463_),
    .A2(_1457_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3899_ (.A1(_1462_),
    .A2(_1455_),
    .B(_1464_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3900_ (.I(_1314_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3901_ (.I(_1150_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3902_ (.A1(_1466_),
    .A2(_1457_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3903_ (.A1(_1465_),
    .A2(_1455_),
    .B(_1467_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3904_ (.I(_1318_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3905_ (.I(_1444_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3906_ (.I(_1155_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3907_ (.I(_1446_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3908_ (.A1(_1470_),
    .A2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3909_ (.A1(_1468_),
    .A2(_1469_),
    .B(_1472_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3910_ (.I(_1324_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3911_ (.I(_1160_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3912_ (.A1(_1474_),
    .A2(_1471_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3913_ (.A1(_1473_),
    .A2(_1469_),
    .B(_1475_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3914_ (.I(_1328_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3915_ (.A1(_1376_),
    .A2(_1471_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3916_ (.A1(_1476_),
    .A2(_1469_),
    .B(_1477_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3917_ (.I(_1165_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3918_ (.A1(_1478_),
    .A2(_1471_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3919_ (.A1(_1379_),
    .A2(_1469_),
    .B(_1479_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3920_ (.I(_1333_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3921_ (.I(_1444_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3922_ (.I(_1170_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3923_ (.I(_1446_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3924_ (.A1(_1482_),
    .A2(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3925_ (.A1(_1480_),
    .A2(_1481_),
    .B(_1484_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3926_ (.I(_1339_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3927_ (.I(_1175_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3928_ (.A1(_1486_),
    .A2(_1483_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3929_ (.A1(_1485_),
    .A2(_1481_),
    .B(_1487_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3930_ (.I(_1343_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3931_ (.I(_1179_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3932_ (.A1(_1489_),
    .A2(_1483_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3933_ (.A1(_1488_),
    .A2(_1481_),
    .B(_1490_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3934_ (.I(_1347_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3935_ (.I(_1183_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3936_ (.A1(_1492_),
    .A2(_1483_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3937_ (.A1(_1491_),
    .A2(_1481_),
    .B(_1493_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3938_ (.A1(_1186_),
    .A2(_1414_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3939_ (.I(_1494_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3940_ (.I(_1495_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3941_ (.I(_1190_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3942_ (.I(_1494_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3943_ (.I(_1498_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3944_ (.A1(_1497_),
    .A2(_1499_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3945_ (.A1(_1442_),
    .A2(_1496_),
    .B(_1500_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3946_ (.I(_1195_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3947_ (.A1(_1501_),
    .A2(_1499_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3948_ (.A1(_1449_),
    .A2(_1496_),
    .B(_1502_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3949_ (.I(_1198_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3950_ (.A1(_1503_),
    .A2(_1499_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3951_ (.A1(_1451_),
    .A2(_1496_),
    .B(_1504_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3952_ (.I(_1201_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3953_ (.A1(_1505_),
    .A2(_1499_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3954_ (.A1(_1453_),
    .A2(_1496_),
    .B(_1506_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3955_ (.I(_1364_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3956_ (.I(_1495_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3957_ (.I(_1498_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3958_ (.A1(_1456_),
    .A2(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3959_ (.A1(_1507_),
    .A2(_1508_),
    .B(_1510_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3960_ (.A1(_1460_),
    .A2(_1509_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3961_ (.A1(_1459_),
    .A2(_1508_),
    .B(_1511_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3962_ (.A1(_1463_),
    .A2(_1509_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3963_ (.A1(_1462_),
    .A2(_1508_),
    .B(_1512_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3964_ (.A1(_1466_),
    .A2(_1509_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3965_ (.A1(_1465_),
    .A2(_1508_),
    .B(_1513_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3966_ (.I(_1495_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3967_ (.I(_1498_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3968_ (.A1(_1470_),
    .A2(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3969_ (.A1(_1468_),
    .A2(_1514_),
    .B(_1516_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3970_ (.A1(_1474_),
    .A2(_1515_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3971_ (.A1(_1473_),
    .A2(_1514_),
    .B(_1517_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3972_ (.I(_1215_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3973_ (.A1(_1518_),
    .A2(_1515_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3974_ (.A1(_1476_),
    .A2(_1514_),
    .B(_1519_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3975_ (.I(_1378_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3976_ (.A1(_1478_),
    .A2(_1515_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3977_ (.A1(_1520_),
    .A2(_1514_),
    .B(_1521_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3978_ (.I(_1495_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3979_ (.I(_1498_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_1482_),
    .A2(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3981_ (.A1(_1480_),
    .A2(_1522_),
    .B(_1524_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3982_ (.A1(_1486_),
    .A2(_1523_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3983_ (.A1(_1485_),
    .A2(_1522_),
    .B(_1525_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3984_ (.A1(_1489_),
    .A2(_1523_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3985_ (.A1(_1488_),
    .A2(_1522_),
    .B(_1526_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3986_ (.A1(_1492_),
    .A2(_1523_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3987_ (.A1(_1491_),
    .A2(_1522_),
    .B(_1527_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3988_ (.I(_0882_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3989_ (.A1(_1528_),
    .A2(_1226_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3990_ (.I(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3991_ (.I(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3992_ (.I(_1529_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3993_ (.I(_1532_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3994_ (.A1(_1497_),
    .A2(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3995_ (.A1(_1442_),
    .A2(_1531_),
    .B(_1534_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3996_ (.A1(_1501_),
    .A2(_1533_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3997_ (.A1(_1449_),
    .A2(_1531_),
    .B(_1535_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3998_ (.A1(_1503_),
    .A2(_1533_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3999_ (.A1(_1451_),
    .A2(_1531_),
    .B(_1536_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4000_ (.A1(_1505_),
    .A2(_1533_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4001_ (.A1(_1453_),
    .A2(_1531_),
    .B(_1537_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4002_ (.I(_1530_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4003_ (.I(_1532_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4004_ (.A1(_1456_),
    .A2(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4005_ (.A1(_1507_),
    .A2(_1538_),
    .B(_1540_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4006_ (.A1(_1460_),
    .A2(_1539_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4007_ (.A1(_1459_),
    .A2(_1538_),
    .B(_1541_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4008_ (.A1(_1463_),
    .A2(_1539_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4009_ (.A1(_1462_),
    .A2(_1538_),
    .B(_1542_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4010_ (.A1(_1466_),
    .A2(_1539_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4011_ (.A1(_1465_),
    .A2(_1538_),
    .B(_1543_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4012_ (.I(_1530_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4013_ (.I(_1532_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4014_ (.A1(_1470_),
    .A2(_1545_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4015_ (.A1(_1468_),
    .A2(_1544_),
    .B(_1546_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4016_ (.A1(_1474_),
    .A2(_1545_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4017_ (.A1(_1473_),
    .A2(_1544_),
    .B(_1547_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4018_ (.A1(_1518_),
    .A2(_1545_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4019_ (.A1(_1476_),
    .A2(_1544_),
    .B(_1548_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4020_ (.A1(_1478_),
    .A2(_1545_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4021_ (.A1(_1520_),
    .A2(_1544_),
    .B(_1549_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4022_ (.I(_1530_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4023_ (.I(_1532_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4024_ (.A1(_1482_),
    .A2(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4025_ (.A1(_1480_),
    .A2(_1550_),
    .B(_1552_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4026_ (.A1(_1486_),
    .A2(_1551_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4027_ (.A1(_1485_),
    .A2(_1550_),
    .B(_1553_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4028_ (.A1(_1489_),
    .A2(_1551_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4029_ (.A1(_1488_),
    .A2(_1550_),
    .B(_1554_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4030_ (.A1(_1492_),
    .A2(_1551_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4031_ (.A1(_1491_),
    .A2(_1550_),
    .B(_1555_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4032_ (.A1(_1528_),
    .A2(_0931_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4033_ (.I(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4034_ (.I(_1557_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4035_ (.I(_1556_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4036_ (.I(_1559_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4037_ (.A1(_1497_),
    .A2(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4038_ (.A1(_1442_),
    .A2(_1558_),
    .B(_1561_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4039_ (.A1(_1501_),
    .A2(_1560_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4040_ (.A1(_1449_),
    .A2(_1558_),
    .B(_1562_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4041_ (.A1(_1503_),
    .A2(_1560_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4042_ (.A1(_1451_),
    .A2(_1558_),
    .B(_1563_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4043_ (.A1(_1505_),
    .A2(_1560_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4044_ (.A1(_1453_),
    .A2(_1558_),
    .B(_1564_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4045_ (.I(_1557_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4046_ (.I(_1559_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4047_ (.A1(_1456_),
    .A2(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4048_ (.A1(_1507_),
    .A2(_1565_),
    .B(_1567_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4049_ (.A1(_1460_),
    .A2(_1566_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4050_ (.A1(_1459_),
    .A2(_1565_),
    .B(_1568_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4051_ (.A1(_1463_),
    .A2(_1566_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4052_ (.A1(_1462_),
    .A2(_1565_),
    .B(_1569_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4053_ (.A1(_1466_),
    .A2(_1566_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4054_ (.A1(_1465_),
    .A2(_1565_),
    .B(_1570_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4055_ (.I(_1557_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4056_ (.I(_1559_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4057_ (.A1(_1470_),
    .A2(_1572_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4058_ (.A1(_1468_),
    .A2(_1571_),
    .B(_1573_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4059_ (.A1(_1474_),
    .A2(_1572_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4060_ (.A1(_1473_),
    .A2(_1571_),
    .B(_1574_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4061_ (.A1(_1518_),
    .A2(_1572_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4062_ (.A1(_1476_),
    .A2(_1571_),
    .B(_1575_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4063_ (.A1(_1478_),
    .A2(_1572_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4064_ (.A1(_1520_),
    .A2(_1571_),
    .B(_1576_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4065_ (.I(_1557_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4066_ (.I(_1559_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4067_ (.A1(_1482_),
    .A2(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4068_ (.A1(_1480_),
    .A2(_1577_),
    .B(_1579_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4069_ (.A1(_1486_),
    .A2(_1578_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4070_ (.A1(_1485_),
    .A2(_1577_),
    .B(_1580_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4071_ (.A1(_1489_),
    .A2(_1578_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4072_ (.A1(_1488_),
    .A2(_1577_),
    .B(_1581_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4073_ (.A1(_1492_),
    .A2(_1578_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4074_ (.A1(_1491_),
    .A2(_1577_),
    .B(_1582_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4075_ (.I(_1284_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4076_ (.A1(_1528_),
    .A2(_1286_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4077_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4078_ (.I(_1585_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4079_ (.I(_1584_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4080_ (.I(_1587_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4081_ (.A1(_1497_),
    .A2(_1588_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4082_ (.A1(_1583_),
    .A2(_1586_),
    .B(_1589_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4083_ (.I(_1293_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4084_ (.A1(_1501_),
    .A2(_1588_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4085_ (.A1(_1590_),
    .A2(_1586_),
    .B(_1591_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4086_ (.I(_1296_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4087_ (.A1(_1503_),
    .A2(_1588_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4088_ (.A1(_1592_),
    .A2(_1586_),
    .B(_1593_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4089_ (.I(_1299_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4090_ (.A1(_1505_),
    .A2(_1588_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4091_ (.A1(_1594_),
    .A2(_1586_),
    .B(_1595_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4092_ (.I(_1585_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4093_ (.I(_1137_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4094_ (.I(_1587_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4095_ (.A1(_1597_),
    .A2(_1598_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4096_ (.A1(_1507_),
    .A2(_1596_),
    .B(_1599_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4097_ (.I(_1306_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4098_ (.I(_1142_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4099_ (.A1(_1601_),
    .A2(_1598_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4100_ (.A1(_1600_),
    .A2(_1596_),
    .B(_1602_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4101_ (.I(_1310_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4102_ (.I(_1146_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4103_ (.A1(_1604_),
    .A2(_1598_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4104_ (.A1(_1603_),
    .A2(_1596_),
    .B(_1605_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4105_ (.I(_1314_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4106_ (.I(_1150_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4107_ (.A1(_1607_),
    .A2(_1598_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4108_ (.A1(_1606_),
    .A2(_1596_),
    .B(_1608_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4109_ (.I(_1318_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4110_ (.I(_1585_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4111_ (.I(_1155_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4112_ (.I(_1587_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4113_ (.A1(_1611_),
    .A2(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4114_ (.A1(_1609_),
    .A2(_1610_),
    .B(_1613_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4115_ (.I(_1324_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4116_ (.I(_1160_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4117_ (.A1(_1615_),
    .A2(_1612_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4118_ (.A1(_1614_),
    .A2(_1610_),
    .B(_1616_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4119_ (.I(_1328_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4120_ (.A1(_1518_),
    .A2(_1612_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4121_ (.A1(_1617_),
    .A2(_1610_),
    .B(_1618_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4122_ (.I(_1165_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4123_ (.A1(_1619_),
    .A2(_1612_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4124_ (.A1(_1520_),
    .A2(_1610_),
    .B(_1620_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4125_ (.I(_1333_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4126_ (.I(_1585_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4127_ (.I(_1170_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4128_ (.I(_1587_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4129_ (.A1(_1623_),
    .A2(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4130_ (.A1(_1621_),
    .A2(_1622_),
    .B(_1625_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4131_ (.I(_1339_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4132_ (.I(_1175_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4133_ (.A1(_1627_),
    .A2(_1624_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4134_ (.A1(_1626_),
    .A2(_1622_),
    .B(_1628_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4135_ (.I(_1343_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4136_ (.I(_1179_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4137_ (.A1(_1630_),
    .A2(_1624_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4138_ (.A1(_1629_),
    .A2(_1622_),
    .B(_1631_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4139_ (.I(_1347_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4140_ (.I(_1183_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4141_ (.A1(_1633_),
    .A2(_1624_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4142_ (.A1(_1632_),
    .A2(_1622_),
    .B(_1634_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4143_ (.A1(_1528_),
    .A2(_1033_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4144_ (.I(_1635_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4145_ (.I(_1636_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4146_ (.I(_1190_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4147_ (.I(_1635_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4148_ (.I(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4149_ (.A1(_1638_),
    .A2(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4150_ (.A1(_1583_),
    .A2(_1637_),
    .B(_1641_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4151_ (.I(_1195_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4152_ (.A1(_1642_),
    .A2(_1640_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4153_ (.A1(_1590_),
    .A2(_1637_),
    .B(_1643_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4154_ (.I(_1198_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(_1644_),
    .A2(_1640_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4156_ (.A1(_1592_),
    .A2(_1637_),
    .B(_1645_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4157_ (.I(_1201_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4158_ (.A1(_1646_),
    .A2(_1640_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4159_ (.A1(_1594_),
    .A2(_1637_),
    .B(_1647_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4160_ (.I(_1364_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4161_ (.I(_1636_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4162_ (.I(_1639_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4163_ (.A1(_1597_),
    .A2(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4164_ (.A1(_1648_),
    .A2(_1649_),
    .B(_1651_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4165_ (.A1(_1601_),
    .A2(_1650_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4166_ (.A1(_1600_),
    .A2(_1649_),
    .B(_1652_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4167_ (.A1(_1604_),
    .A2(_1650_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4168_ (.A1(_1603_),
    .A2(_1649_),
    .B(_1653_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4169_ (.A1(_1607_),
    .A2(_1650_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4170_ (.A1(_1606_),
    .A2(_1649_),
    .B(_1654_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4171_ (.I(_1636_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4172_ (.I(_1639_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4173_ (.A1(_1611_),
    .A2(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4174_ (.A1(_1609_),
    .A2(_1655_),
    .B(_1657_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4175_ (.A1(_1615_),
    .A2(_1656_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4176_ (.A1(_1614_),
    .A2(_1655_),
    .B(_1658_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4177_ (.I(_1215_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4178_ (.A1(_1659_),
    .A2(_1656_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4179_ (.A1(_1617_),
    .A2(_1655_),
    .B(_1660_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4180_ (.I(_1378_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4181_ (.A1(_1619_),
    .A2(_1656_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4182_ (.A1(_1661_),
    .A2(_1655_),
    .B(_1662_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4183_ (.I(_1636_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4184_ (.I(_1639_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4185_ (.A1(_1623_),
    .A2(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4186_ (.A1(_1621_),
    .A2(_1663_),
    .B(_1665_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4187_ (.A1(_1627_),
    .A2(_1664_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4188_ (.A1(_1626_),
    .A2(_1663_),
    .B(_1666_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4189_ (.A1(_1630_),
    .A2(_1664_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4190_ (.A1(_1629_),
    .A2(_1663_),
    .B(_1667_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(_1633_),
    .A2(_1664_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4192_ (.A1(_1632_),
    .A2(_1663_),
    .B(_1668_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4193_ (.A1(_0883_),
    .A2(_1068_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4194_ (.I(_1669_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4195_ (.I(_1670_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4196_ (.I(_1669_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4197_ (.I(_1672_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4198_ (.A1(_1638_),
    .A2(_1673_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4199_ (.A1(_1583_),
    .A2(_1671_),
    .B(_1674_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4200_ (.A1(_1642_),
    .A2(_1673_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4201_ (.A1(_1590_),
    .A2(_1671_),
    .B(_1675_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4202_ (.A1(_1644_),
    .A2(_1673_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4203_ (.A1(_1592_),
    .A2(_1671_),
    .B(_1676_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4204_ (.A1(_1646_),
    .A2(_1673_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4205_ (.A1(_1594_),
    .A2(_1671_),
    .B(_1677_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4206_ (.I(_1670_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4207_ (.I(_1672_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4208_ (.A1(_1597_),
    .A2(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4209_ (.A1(_1648_),
    .A2(_1678_),
    .B(_1680_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4210_ (.A1(_1601_),
    .A2(_1679_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4211_ (.A1(_1600_),
    .A2(_1678_),
    .B(_1681_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4212_ (.A1(_1604_),
    .A2(_1679_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4213_ (.A1(_1603_),
    .A2(_1678_),
    .B(_1682_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4214_ (.A1(_1607_),
    .A2(_1679_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4215_ (.A1(_1606_),
    .A2(_1678_),
    .B(_1683_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4216_ (.I(_1670_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4217_ (.I(_1672_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4218_ (.A1(_1611_),
    .A2(_1685_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4219_ (.A1(_1609_),
    .A2(_1684_),
    .B(_1686_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4220_ (.A1(_1615_),
    .A2(_1685_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4221_ (.A1(_1614_),
    .A2(_1684_),
    .B(_1687_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4222_ (.A1(_1659_),
    .A2(_1685_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4223_ (.A1(_1617_),
    .A2(_1684_),
    .B(_1688_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4224_ (.A1(_1619_),
    .A2(_1685_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4225_ (.A1(_1661_),
    .A2(_1684_),
    .B(_1689_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4226_ (.I(_1670_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4227_ (.I(_1672_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4228_ (.A1(_1623_),
    .A2(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4229_ (.A1(_1621_),
    .A2(_1690_),
    .B(_1692_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4230_ (.A1(_1627_),
    .A2(_1691_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4231_ (.A1(_1626_),
    .A2(_1690_),
    .B(_1693_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4232_ (.A1(_1630_),
    .A2(_1691_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4233_ (.A1(_1629_),
    .A2(_1690_),
    .B(_1694_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4234_ (.A1(_1633_),
    .A2(_1691_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4235_ (.A1(_1632_),
    .A2(_1690_),
    .B(_1695_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4236_ (.A1(_0883_),
    .A2(_0964_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4237_ (.I(_1696_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4238_ (.I(_1697_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4239_ (.I(_1696_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4240_ (.I(_1699_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4241_ (.A1(_1638_),
    .A2(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4242_ (.A1(_1583_),
    .A2(_1698_),
    .B(_1701_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4243_ (.A1(_1642_),
    .A2(_1700_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4244_ (.A1(_1590_),
    .A2(_1698_),
    .B(_1702_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4245_ (.A1(_1644_),
    .A2(_1700_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4246_ (.A1(_1592_),
    .A2(_1698_),
    .B(_1703_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4247_ (.A1(_1646_),
    .A2(_1700_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4248_ (.A1(_1594_),
    .A2(_1698_),
    .B(_1704_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4249_ (.I(_1697_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4250_ (.I(_1699_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4251_ (.A1(_1597_),
    .A2(_1706_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4252_ (.A1(_1648_),
    .A2(_1705_),
    .B(_1707_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4253_ (.A1(_1601_),
    .A2(_1706_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4254_ (.A1(_1600_),
    .A2(_1705_),
    .B(_1708_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4255_ (.A1(_1604_),
    .A2(_1706_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4256_ (.A1(_1603_),
    .A2(_1705_),
    .B(_1709_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4257_ (.A1(_1607_),
    .A2(_1706_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4258_ (.A1(_1606_),
    .A2(_1705_),
    .B(_1710_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4259_ (.I(_1697_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4260_ (.I(_1699_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4261_ (.A1(_1611_),
    .A2(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4262_ (.A1(_1609_),
    .A2(_1711_),
    .B(_1713_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4263_ (.A1(_1615_),
    .A2(_1712_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4264_ (.A1(_1614_),
    .A2(_1711_),
    .B(_1714_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4265_ (.A1(_1659_),
    .A2(_1712_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4266_ (.A1(_1617_),
    .A2(_1711_),
    .B(_1715_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4267_ (.A1(_1619_),
    .A2(_1712_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4268_ (.A1(_1661_),
    .A2(_1711_),
    .B(_1716_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4269_ (.I(_1697_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4270_ (.I(_1699_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4271_ (.A1(_1623_),
    .A2(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4272_ (.A1(_1621_),
    .A2(_1717_),
    .B(_1719_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4273_ (.A1(_1627_),
    .A2(_1718_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4274_ (.A1(_1626_),
    .A2(_1717_),
    .B(_1720_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4275_ (.A1(_1630_),
    .A2(_1718_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4276_ (.A1(_1629_),
    .A2(_1717_),
    .B(_1721_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4277_ (.A1(_1633_),
    .A2(_1718_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4278_ (.A1(_1632_),
    .A2(_1717_),
    .B(_1722_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4279_ (.I(_1284_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4280_ (.I(_0965_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4281_ (.A1(_1724_),
    .A2(_1186_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4282_ (.I(_1725_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4283_ (.I(_1726_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4284_ (.I(_1725_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4285_ (.I(_1728_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4286_ (.A1(_1638_),
    .A2(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4287_ (.A1(_1723_),
    .A2(_1727_),
    .B(_1730_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4288_ (.I(_1293_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4289_ (.A1(_1642_),
    .A2(_1729_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4290_ (.A1(_1731_),
    .A2(_1727_),
    .B(_1732_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4291_ (.I(_1296_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_1644_),
    .A2(_1729_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4293_ (.A1(_1733_),
    .A2(_1727_),
    .B(_1734_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4294_ (.I(_1299_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4295_ (.A1(_1646_),
    .A2(_1729_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4296_ (.A1(_1735_),
    .A2(_1727_),
    .B(_1736_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4297_ (.I(_1726_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4298_ (.I(net28),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4299_ (.I(_1728_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4300_ (.A1(_1738_),
    .A2(_1739_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4301_ (.A1(_1648_),
    .A2(_1737_),
    .B(_1740_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4302_ (.I(_1306_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4303_ (.I(net29),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4304_ (.A1(_1742_),
    .A2(_1739_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4305_ (.A1(_1741_),
    .A2(_1737_),
    .B(_1743_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4306_ (.I(_1310_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4307_ (.I(net30),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4308_ (.A1(_1745_),
    .A2(_1739_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4309_ (.A1(_1744_),
    .A2(_1737_),
    .B(_1746_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4310_ (.I(_1314_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4311_ (.I(net31),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4312_ (.A1(_1748_),
    .A2(_1739_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4313_ (.A1(_1747_),
    .A2(_1737_),
    .B(_1749_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4314_ (.I(_1318_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4315_ (.I(_1726_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4316_ (.I(net32),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4317_ (.I(_1728_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4318_ (.A1(_1752_),
    .A2(_1753_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4319_ (.A1(_1750_),
    .A2(_1751_),
    .B(_1754_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4320_ (.I(_1324_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4321_ (.I(net33),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4322_ (.A1(_1756_),
    .A2(_1753_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4323_ (.A1(_1755_),
    .A2(_1751_),
    .B(_1757_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4324_ (.I(_1328_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4325_ (.A1(_1659_),
    .A2(_1753_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4326_ (.A1(_1758_),
    .A2(_1751_),
    .B(_1759_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4327_ (.I(net20),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4328_ (.A1(_1760_),
    .A2(_1753_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4329_ (.A1(_1661_),
    .A2(_1751_),
    .B(_1761_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4330_ (.I(_1333_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4331_ (.I(_1726_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4332_ (.I(net21),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4333_ (.I(_1728_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4334_ (.A1(_1764_),
    .A2(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4335_ (.A1(_1762_),
    .A2(_1763_),
    .B(_1766_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4336_ (.I(_1339_),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4337_ (.I(net22),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4338_ (.A1(_1768_),
    .A2(_1765_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4339_ (.A1(_1767_),
    .A2(_1763_),
    .B(_1769_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4340_ (.I(_1343_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4341_ (.I(net23),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4342_ (.A1(_1771_),
    .A2(_1765_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4343_ (.A1(_1770_),
    .A2(_1763_),
    .B(_1772_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4344_ (.I(_1347_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4345_ (.I(net24),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4346_ (.A1(_1774_),
    .A2(_1765_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4347_ (.A1(_1773_),
    .A2(_1763_),
    .B(_1775_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4348_ (.A1(_0883_),
    .A2(_1186_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4349_ (.I(_1776_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4350_ (.I(_1777_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4351_ (.I(net18),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4352_ (.I(_1776_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4353_ (.I(_1780_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4354_ (.A1(_1779_),
    .A2(_1781_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4355_ (.A1(_1723_),
    .A2(_1778_),
    .B(_1782_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4356_ (.I(net25),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4357_ (.A1(_1783_),
    .A2(_1781_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4358_ (.A1(_1731_),
    .A2(_1778_),
    .B(_1784_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4359_ (.I(net26),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4360_ (.A1(_1785_),
    .A2(_1781_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4361_ (.A1(_1733_),
    .A2(_1778_),
    .B(_1786_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4362_ (.I(net27),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4363_ (.A1(_1787_),
    .A2(_1781_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4364_ (.A1(_1735_),
    .A2(_1778_),
    .B(_1788_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4365_ (.I(_1364_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4366_ (.I(_1777_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4367_ (.I(_1780_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4368_ (.A1(_1738_),
    .A2(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4369_ (.A1(_1789_),
    .A2(_1790_),
    .B(_1792_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4370_ (.A1(_1742_),
    .A2(_1791_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4371_ (.A1(_1741_),
    .A2(_1790_),
    .B(_1793_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4372_ (.A1(_1745_),
    .A2(_1791_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4373_ (.A1(_1744_),
    .A2(_1790_),
    .B(_1794_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4374_ (.A1(_1748_),
    .A2(_1791_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4375_ (.A1(_1747_),
    .A2(_1790_),
    .B(_1795_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4376_ (.I(_1777_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4377_ (.I(_1780_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4378_ (.A1(_1752_),
    .A2(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4379_ (.A1(_1750_),
    .A2(_1796_),
    .B(_1798_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4380_ (.A1(_1756_),
    .A2(_1797_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4381_ (.A1(_1755_),
    .A2(_1796_),
    .B(_1799_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4382_ (.I(net19),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4383_ (.A1(_1800_),
    .A2(_1797_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4384_ (.A1(_1758_),
    .A2(_1796_),
    .B(_1801_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4385_ (.I(_1378_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4386_ (.A1(_1760_),
    .A2(_1797_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4387_ (.A1(_1802_),
    .A2(_1796_),
    .B(_1803_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4388_ (.I(_1777_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4389_ (.I(_1780_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4390_ (.A1(_1764_),
    .A2(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4391_ (.A1(_1762_),
    .A2(_1804_),
    .B(_1806_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4392_ (.A1(_1768_),
    .A2(_1805_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4393_ (.A1(_1767_),
    .A2(_1804_),
    .B(_1807_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4394_ (.A1(_1771_),
    .A2(_1805_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4395_ (.A1(_1770_),
    .A2(_1804_),
    .B(_1808_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4396_ (.A1(_1774_),
    .A2(_1805_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4397_ (.A1(_1773_),
    .A2(_1804_),
    .B(_1809_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4398_ (.A1(_1724_),
    .A2(_1226_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4399_ (.I(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4400_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4401_ (.I(_1810_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4402_ (.I(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4403_ (.A1(_1779_),
    .A2(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4404_ (.A1(_1723_),
    .A2(_1812_),
    .B(_1815_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4405_ (.A1(_1783_),
    .A2(_1814_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4406_ (.A1(_1731_),
    .A2(_1812_),
    .B(_1816_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4407_ (.A1(_1785_),
    .A2(_1814_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4408_ (.A1(_1733_),
    .A2(_1812_),
    .B(_1817_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4409_ (.A1(_1787_),
    .A2(_1814_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4410_ (.A1(_1735_),
    .A2(_1812_),
    .B(_1818_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4411_ (.I(_1811_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4412_ (.I(_1813_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4413_ (.A1(_1738_),
    .A2(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4414_ (.A1(_1789_),
    .A2(_1819_),
    .B(_1821_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4415_ (.A1(_1742_),
    .A2(_1820_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4416_ (.A1(_1741_),
    .A2(_1819_),
    .B(_1822_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4417_ (.A1(_1745_),
    .A2(_1820_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4418_ (.A1(_1744_),
    .A2(_1819_),
    .B(_1823_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4419_ (.A1(_1748_),
    .A2(_1820_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4420_ (.A1(_1747_),
    .A2(_1819_),
    .B(_1824_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4421_ (.I(_1811_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4422_ (.I(_1813_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4423_ (.A1(_1752_),
    .A2(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4424_ (.A1(_1750_),
    .A2(_1825_),
    .B(_1827_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4425_ (.A1(_1756_),
    .A2(_1826_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4426_ (.A1(_1755_),
    .A2(_1825_),
    .B(_1828_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4427_ (.A1(_1800_),
    .A2(_1826_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4428_ (.A1(_1758_),
    .A2(_1825_),
    .B(_1829_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4429_ (.A1(_1760_),
    .A2(_1826_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4430_ (.A1(_1802_),
    .A2(_1825_),
    .B(_1830_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4431_ (.I(_1811_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4432_ (.I(_1813_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4433_ (.A1(_1764_),
    .A2(_1832_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4434_ (.A1(_1762_),
    .A2(_1831_),
    .B(_1833_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4435_ (.A1(_1768_),
    .A2(_1832_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4436_ (.A1(_1767_),
    .A2(_1831_),
    .B(_1834_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4437_ (.A1(_1771_),
    .A2(_1832_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4438_ (.A1(_1770_),
    .A2(_1831_),
    .B(_1835_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4439_ (.A1(_1774_),
    .A2(_1832_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4440_ (.A1(_1773_),
    .A2(_1831_),
    .B(_1836_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(_0931_),
    .A2(_0966_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4442_ (.I(_1837_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4443_ (.I(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4444_ (.I(_1837_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4445_ (.I(_1840_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4446_ (.A1(_1779_),
    .A2(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4447_ (.A1(_1723_),
    .A2(_1839_),
    .B(_1842_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4448_ (.A1(_1783_),
    .A2(_1841_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4449_ (.A1(_1731_),
    .A2(_1839_),
    .B(_1843_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4450_ (.A1(_1785_),
    .A2(_1841_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4451_ (.A1(_1733_),
    .A2(_1839_),
    .B(_1844_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4452_ (.A1(_1787_),
    .A2(_1841_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4453_ (.A1(_1735_),
    .A2(_1839_),
    .B(_1845_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4454_ (.I(_1838_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4455_ (.I(_1840_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4456_ (.A1(_1738_),
    .A2(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4457_ (.A1(_1789_),
    .A2(_1846_),
    .B(_1848_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4458_ (.A1(_1742_),
    .A2(_1847_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4459_ (.A1(_1741_),
    .A2(_1846_),
    .B(_1849_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4460_ (.A1(_1745_),
    .A2(_1847_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4461_ (.A1(_1744_),
    .A2(_1846_),
    .B(_1850_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4462_ (.A1(_1748_),
    .A2(_1847_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4463_ (.A1(_1747_),
    .A2(_1846_),
    .B(_1851_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4464_ (.I(_1838_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4465_ (.I(_1840_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4466_ (.A1(_1752_),
    .A2(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4467_ (.A1(_1750_),
    .A2(_1852_),
    .B(_1854_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4468_ (.A1(_1756_),
    .A2(_1853_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4469_ (.A1(_1755_),
    .A2(_1852_),
    .B(_1855_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4470_ (.A1(_1800_),
    .A2(_1853_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4471_ (.A1(_1758_),
    .A2(_1852_),
    .B(_1856_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4472_ (.A1(_1760_),
    .A2(_1853_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4473_ (.A1(_1802_),
    .A2(_1852_),
    .B(_1857_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4474_ (.I(_1838_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4475_ (.I(_1840_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4476_ (.A1(_1764_),
    .A2(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4477_ (.A1(_1762_),
    .A2(_1858_),
    .B(_1860_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4478_ (.A1(_1768_),
    .A2(_1859_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4479_ (.A1(_1767_),
    .A2(_1858_),
    .B(_1861_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4480_ (.A1(_1771_),
    .A2(_1859_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4481_ (.A1(_1770_),
    .A2(_1858_),
    .B(_1862_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4482_ (.A1(_1774_),
    .A2(_1859_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4483_ (.A1(_1773_),
    .A2(_1858_),
    .B(_1863_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4484_ (.I(_2145_),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4485_ (.A1(_1724_),
    .A2(_1286_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4486_ (.I(_1865_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4487_ (.I(_1866_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4488_ (.I(_1865_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4489_ (.I(_1868_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4490_ (.A1(_1779_),
    .A2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4491_ (.A1(_1864_),
    .A2(_1867_),
    .B(_1870_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4492_ (.I(_2171_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4493_ (.A1(_1783_),
    .A2(_1869_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4494_ (.A1(_1871_),
    .A2(_1867_),
    .B(_1872_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4495_ (.I(_2189_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4496_ (.A1(_1785_),
    .A2(_1869_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4497_ (.A1(_1873_),
    .A2(_1867_),
    .B(_1874_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4498_ (.I(_2211_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4499_ (.A1(_1787_),
    .A2(_1869_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4500_ (.A1(_1875_),
    .A2(_1867_),
    .B(_1876_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4501_ (.I(_1866_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4502_ (.I(net28),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4503_ (.I(_1868_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4504_ (.A1(_1878_),
    .A2(_1879_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4505_ (.A1(_1789_),
    .A2(_1877_),
    .B(_1880_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4506_ (.I(_2256_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4507_ (.I(net29),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4508_ (.A1(_1882_),
    .A2(_1879_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4509_ (.A1(_1881_),
    .A2(_1877_),
    .B(_1883_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4510_ (.I(_2277_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4511_ (.I(net30),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4512_ (.A1(_1885_),
    .A2(_1879_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4513_ (.A1(_1884_),
    .A2(_1877_),
    .B(_1886_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4514_ (.I(_2297_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4515_ (.I(net31),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4516_ (.A1(_1888_),
    .A2(_1879_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4517_ (.A1(_1887_),
    .A2(_1877_),
    .B(_1889_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4518_ (.I(_2321_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4519_ (.I(_1866_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4520_ (.I(net32),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4521_ (.I(_1868_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4522_ (.A1(_1892_),
    .A2(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4523_ (.A1(_1890_),
    .A2(_1891_),
    .B(_1894_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4524_ (.I(_2335_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4525_ (.I(net33),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4526_ (.A1(_1896_),
    .A2(_1893_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4527_ (.A1(_1895_),
    .A2(_1891_),
    .B(_1897_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4528_ (.I(_2354_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4529_ (.A1(_1800_),
    .A2(_1893_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4530_ (.A1(_1898_),
    .A2(_1891_),
    .B(_1899_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4531_ (.I(net20),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4532_ (.A1(_1900_),
    .A2(_1893_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4533_ (.A1(_1802_),
    .A2(_1891_),
    .B(_1901_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4534_ (.I(_0571_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4535_ (.I(_1866_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4536_ (.I(net21),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4537_ (.I(_1868_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4538_ (.A1(_1904_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4539_ (.A1(_1902_),
    .A2(_1903_),
    .B(_1906_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4540_ (.I(_0591_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4541_ (.I(net22),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4542_ (.A1(_1908_),
    .A2(_1905_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4543_ (.A1(_1907_),
    .A2(_1903_),
    .B(_1909_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4544_ (.I(_0603_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4545_ (.I(net23),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4546_ (.A1(_1911_),
    .A2(_1905_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4547_ (.A1(_1910_),
    .A2(_1903_),
    .B(_1912_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_0614_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4549_ (.I(net24),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4550_ (.A1(_1914_),
    .A2(_1905_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4551_ (.A1(_1913_),
    .A2(_1903_),
    .B(_1915_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4552_ (.A1(_1724_),
    .A2(_1033_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4553_ (.I(_1916_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4555_ (.I(net18),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4556_ (.I(_1916_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4557_ (.I(_1920_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4558_ (.A1(_1919_),
    .A2(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4559_ (.A1(_1864_),
    .A2(_1918_),
    .B(_1922_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4560_ (.I(net25),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4561_ (.A1(_1923_),
    .A2(_1921_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4562_ (.A1(_1871_),
    .A2(_1918_),
    .B(_1924_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4563_ (.I(net26),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4564_ (.A1(_1925_),
    .A2(_1921_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4565_ (.A1(_1873_),
    .A2(_1918_),
    .B(_1926_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4566_ (.I(net27),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4567_ (.A1(_1927_),
    .A2(_1921_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4568_ (.A1(_1875_),
    .A2(_1918_),
    .B(_1928_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4569_ (.I(_2232_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4570_ (.I(_1917_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4571_ (.I(_1920_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4572_ (.A1(_1878_),
    .A2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4573_ (.A1(_1929_),
    .A2(_1930_),
    .B(_1932_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4574_ (.A1(_1882_),
    .A2(_1931_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4575_ (.A1(_1881_),
    .A2(_1930_),
    .B(_1933_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4576_ (.A1(_1885_),
    .A2(_1931_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4577_ (.A1(_1884_),
    .A2(_1930_),
    .B(_1934_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4578_ (.A1(_1888_),
    .A2(_1931_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4579_ (.A1(_1887_),
    .A2(_1930_),
    .B(_1935_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_1917_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(_1920_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4582_ (.A1(_1892_),
    .A2(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4583_ (.A1(_1890_),
    .A2(_1936_),
    .B(_1938_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_1896_),
    .A2(_1937_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4585_ (.A1(_1895_),
    .A2(_1936_),
    .B(_1939_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4586_ (.I(net19),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4587_ (.A1(_1940_),
    .A2(_1937_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4588_ (.A1(_1898_),
    .A2(_1936_),
    .B(_1941_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4589_ (.I(_2370_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4590_ (.A1(_1900_),
    .A2(_1937_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4591_ (.A1(_1942_),
    .A2(_1936_),
    .B(_1943_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4592_ (.I(_1917_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4593_ (.I(_1920_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4594_ (.A1(_1904_),
    .A2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4595_ (.A1(_1902_),
    .A2(_1944_),
    .B(_1946_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4596_ (.A1(_1908_),
    .A2(_1945_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4597_ (.A1(_1907_),
    .A2(_1944_),
    .B(_1947_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4598_ (.A1(_1911_),
    .A2(_1945_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4599_ (.A1(_1910_),
    .A2(_1944_),
    .B(_1948_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4600_ (.A1(_1914_),
    .A2(_1945_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4601_ (.A1(_1913_),
    .A2(_1944_),
    .B(_1949_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4602_ (.A1(_0966_),
    .A2(_1068_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4603_ (.I(_1950_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4604_ (.I(_1951_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4605_ (.I(_1950_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4606_ (.I(_1953_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4607_ (.A1(_1919_),
    .A2(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4608_ (.A1(_1864_),
    .A2(_1952_),
    .B(_1955_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4609_ (.A1(_1923_),
    .A2(_1954_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4610_ (.A1(_1871_),
    .A2(_1952_),
    .B(_1956_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4611_ (.A1(_1925_),
    .A2(_1954_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4612_ (.A1(_1873_),
    .A2(_1952_),
    .B(_1957_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4613_ (.A1(_1927_),
    .A2(_1954_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4614_ (.A1(_1875_),
    .A2(_1952_),
    .B(_1958_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4615_ (.I(_1951_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4616_ (.I(_1953_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4617_ (.A1(_1878_),
    .A2(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4618_ (.A1(_1929_),
    .A2(_1959_),
    .B(_1961_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4619_ (.A1(_1882_),
    .A2(_1960_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4620_ (.A1(_1881_),
    .A2(_1959_),
    .B(_1962_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4621_ (.A1(_1885_),
    .A2(_1960_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4622_ (.A1(_1884_),
    .A2(_1959_),
    .B(_1963_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4623_ (.A1(_1888_),
    .A2(_1960_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4624_ (.A1(_1887_),
    .A2(_1959_),
    .B(_1964_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4625_ (.I(_1951_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4626_ (.I(_1953_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4627_ (.A1(_1892_),
    .A2(_1966_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4628_ (.A1(_1890_),
    .A2(_1965_),
    .B(_1967_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4629_ (.A1(_1896_),
    .A2(_1966_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4630_ (.A1(_1895_),
    .A2(_1965_),
    .B(_1968_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4631_ (.A1(_1940_),
    .A2(_1966_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4632_ (.A1(_1898_),
    .A2(_1965_),
    .B(_1969_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4633_ (.A1(_1900_),
    .A2(_1966_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4634_ (.A1(_1942_),
    .A2(_1965_),
    .B(_1970_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4635_ (.I(_1951_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4636_ (.I(_1953_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4637_ (.A1(_1904_),
    .A2(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4638_ (.A1(_1902_),
    .A2(_1971_),
    .B(_1973_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4639_ (.A1(_1908_),
    .A2(_1972_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4640_ (.A1(_1907_),
    .A2(_1971_),
    .B(_1974_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4641_ (.A1(_1911_),
    .A2(_1972_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4642_ (.A1(_1910_),
    .A2(_1971_),
    .B(_1975_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4643_ (.A1(_1914_),
    .A2(_1972_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4644_ (.A1(_1913_),
    .A2(_1971_),
    .B(_1976_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4645_ (.A1(_0933_),
    .A2(_1226_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4646_ (.I(_1977_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4647_ (.I(_1978_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4648_ (.I(_1977_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4649_ (.I(_1980_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4650_ (.A1(_1919_),
    .A2(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4651_ (.A1(_1864_),
    .A2(_1979_),
    .B(_1982_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4652_ (.A1(_1923_),
    .A2(_1981_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4653_ (.A1(_1871_),
    .A2(_1979_),
    .B(_1983_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4654_ (.A1(_1925_),
    .A2(_1981_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4655_ (.A1(_1873_),
    .A2(_1979_),
    .B(_1984_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4656_ (.A1(_1927_),
    .A2(_1981_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4657_ (.A1(_1875_),
    .A2(_1979_),
    .B(_1985_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4658_ (.I(_1978_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4659_ (.I(_1980_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4660_ (.A1(_1878_),
    .A2(_1987_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4661_ (.A1(_1929_),
    .A2(_1986_),
    .B(_1988_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_1882_),
    .A2(_1987_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4663_ (.A1(_1881_),
    .A2(_1986_),
    .B(_1989_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4664_ (.A1(_1885_),
    .A2(_1987_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4665_ (.A1(_1884_),
    .A2(_1986_),
    .B(_1990_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4666_ (.A1(_1888_),
    .A2(_1987_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4667_ (.A1(_1887_),
    .A2(_1986_),
    .B(_1991_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4668_ (.I(_1978_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4669_ (.I(_1980_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4670_ (.A1(_1892_),
    .A2(_1993_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4671_ (.A1(_1890_),
    .A2(_1992_),
    .B(_1994_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4672_ (.A1(_1896_),
    .A2(_1993_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4673_ (.A1(_1895_),
    .A2(_1992_),
    .B(_1995_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4674_ (.A1(_1940_),
    .A2(_1993_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4675_ (.A1(_1898_),
    .A2(_1992_),
    .B(_1996_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4676_ (.A1(_1900_),
    .A2(_1993_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4677_ (.A1(_1942_),
    .A2(_1992_),
    .B(_1997_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4678_ (.I(_1978_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4679_ (.I(_1980_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4680_ (.A1(_1904_),
    .A2(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4681_ (.A1(_1902_),
    .A2(_1998_),
    .B(_2000_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4682_ (.A1(_1908_),
    .A2(_1999_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4683_ (.A1(_1907_),
    .A2(_1998_),
    .B(_2001_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4684_ (.A1(_1911_),
    .A2(_1999_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4685_ (.A1(_1910_),
    .A2(_1998_),
    .B(_2002_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4686_ (.A1(_1914_),
    .A2(_1999_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4687_ (.A1(_1913_),
    .A2(_1998_),
    .B(_2003_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4688_ (.A1(_0933_),
    .A2(_1286_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4689_ (.I(_2004_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4690_ (.I(_2005_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4691_ (.I(_2004_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4692_ (.I(_2007_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4693_ (.A1(_1919_),
    .A2(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4694_ (.A1(_0961_),
    .A2(_2006_),
    .B(_2009_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4695_ (.A1(_1923_),
    .A2(_2008_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4696_ (.A1(_0973_),
    .A2(_2006_),
    .B(_2010_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4697_ (.A1(_1925_),
    .A2(_2008_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4698_ (.A1(_0976_),
    .A2(_2006_),
    .B(_2011_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4699_ (.A1(_1927_),
    .A2(_2008_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4700_ (.A1(_0979_),
    .A2(_2006_),
    .B(_2012_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4701_ (.I(_2005_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4702_ (.I(_2007_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4703_ (.A1(_0797_),
    .A2(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4704_ (.A1(_1929_),
    .A2(_2013_),
    .B(_2015_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4705_ (.A1(_0801_),
    .A2(_2014_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4706_ (.A1(_0986_),
    .A2(_2013_),
    .B(_2016_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4707_ (.A1(_0804_),
    .A2(_2014_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4708_ (.A1(_0990_),
    .A2(_2013_),
    .B(_2017_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4709_ (.A1(_0807_),
    .A2(_2014_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4710_ (.A1(_0994_),
    .A2(_2013_),
    .B(_2018_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4711_ (.I(_2005_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4712_ (.I(_2007_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4713_ (.A1(_0811_),
    .A2(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4714_ (.A1(_0998_),
    .A2(_2019_),
    .B(_2021_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4715_ (.A1(_0815_),
    .A2(_2020_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4716_ (.A1(_1004_),
    .A2(_2019_),
    .B(_2022_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4717_ (.A1(_1940_),
    .A2(_2020_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4718_ (.A1(_1008_),
    .A2(_2019_),
    .B(_2023_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4719_ (.A1(_0823_),
    .A2(_2020_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4720_ (.A1(_1942_),
    .A2(_2019_),
    .B(_2024_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4721_ (.I(_2005_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4722_ (.I(_2007_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4723_ (.A1(_0827_),
    .A2(_2026_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4724_ (.A1(_1013_),
    .A2(_2025_),
    .B(_2027_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4725_ (.A1(_0831_),
    .A2(_2026_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4726_ (.A1(_1019_),
    .A2(_2025_),
    .B(_2028_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4727_ (.A1(_0834_),
    .A2(_2026_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4728_ (.A1(_1023_),
    .A2(_2025_),
    .B(_2029_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4729_ (.A1(_0837_),
    .A2(_2026_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4730_ (.A1(_1027_),
    .A2(_2025_),
    .B(_2030_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4731_ (.A1(_1068_),
    .A2(_1414_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4732_ (.I(_2031_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4733_ (.I(_2032_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4734_ (.I(_2031_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4735_ (.I(_2034_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4736_ (.A1(_0780_),
    .A2(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4737_ (.A1(_0961_),
    .A2(_2033_),
    .B(_2036_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(_0785_),
    .A2(_2035_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4739_ (.A1(_0973_),
    .A2(_2033_),
    .B(_2037_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4740_ (.A1(_0788_),
    .A2(_2035_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4741_ (.A1(_0976_),
    .A2(_2033_),
    .B(_2038_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4742_ (.A1(_0791_),
    .A2(_2035_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4743_ (.A1(_0979_),
    .A2(_2033_),
    .B(_2039_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4744_ (.I(_2032_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4745_ (.I(_2034_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4746_ (.A1(_0797_),
    .A2(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4747_ (.A1(_0794_),
    .A2(_2040_),
    .B(_2042_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4748_ (.A1(_0801_),
    .A2(_2041_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4749_ (.A1(_0986_),
    .A2(_2040_),
    .B(_2043_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4750_ (.A1(_0804_),
    .A2(_2041_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4751_ (.A1(_0990_),
    .A2(_2040_),
    .B(_2044_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4752_ (.A1(_0807_),
    .A2(_2041_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4753_ (.A1(_0994_),
    .A2(_2040_),
    .B(_2045_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4754_ (.I(_2032_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4755_ (.I(_2034_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4756_ (.A1(_0811_),
    .A2(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4757_ (.A1(_0998_),
    .A2(_2046_),
    .B(_2048_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4758_ (.A1(_0815_),
    .A2(_2047_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4759_ (.A1(_1004_),
    .A2(_2046_),
    .B(_2049_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4760_ (.A1(_0818_),
    .A2(_2047_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4761_ (.A1(_1008_),
    .A2(_2046_),
    .B(_2050_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4762_ (.A1(_0823_),
    .A2(_2047_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4763_ (.A1(_0821_),
    .A2(_2046_),
    .B(_2051_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4764_ (.I(_2032_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4765_ (.I(_2034_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4766_ (.A1(_0827_),
    .A2(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4767_ (.A1(_1013_),
    .A2(_2052_),
    .B(_2054_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4768_ (.A1(_0831_),
    .A2(_2053_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4769_ (.A1(_1019_),
    .A2(_2052_),
    .B(_2055_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4770_ (.A1(_0834_),
    .A2(_2053_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4771_ (.A1(_1023_),
    .A2(_2052_),
    .B(_2056_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4772_ (.A1(_0837_),
    .A2(_2053_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4773_ (.A1(_1027_),
    .A2(_2052_),
    .B(_2057_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4774_ (.I(net47),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4775_ (.A1(_2058_),
    .A2(_0731_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4776_ (.A1(_2145_),
    .A2(_0752_),
    .B1(_0713_),
    .B2(_2119_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4777_ (.A1(net35),
    .A2(_2059_),
    .A3(_2060_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4778_ (.A1(_0718_),
    .A2(_2061_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4779_ (.I(_2062_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4780_ (.I(net51),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4781_ (.A1(_2058_),
    .A2(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4782_ (.A1(_2171_),
    .A2(_0753_),
    .B1(_0732_),
    .B2(_2064_),
    .C(_0708_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4783_ (.A1(_2084_),
    .A2(_0667_),
    .B(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4784_ (.A1(_2063_),
    .A2(_0730_),
    .B(_2066_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4785_ (.I(net52),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4786_ (.A1(_2058_),
    .A2(net51),
    .A3(net52),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4787_ (.A1(_2058_),
    .A2(net51),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4788_ (.A1(_2067_),
    .A2(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4789_ (.A1(_2068_),
    .A2(_2070_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4790_ (.A1(_2189_),
    .A2(_0753_),
    .B1(_0732_),
    .B2(_2071_),
    .C(_0708_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4791_ (.A1(_0688_),
    .A2(_0667_),
    .B(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4792_ (.A1(_2067_),
    .A2(_0730_),
    .B(_2073_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4793_ (.A1(_2211_),
    .A2(_0753_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4794_ (.I(net53),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4795_ (.A1(_2075_),
    .A2(_2068_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4796_ (.A1(\Control_unit2.instr_stage2[3] ),
    .A2(_0747_),
    .B1(_0713_),
    .B2(_2076_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4797_ (.A1(_0709_),
    .A2(_2074_),
    .A3(_2077_),
    .B1(_0749_),
    .B2(_2075_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4798_ (.D(_0000_),
    .RN(net34),
    .CLK(clknet_leaf_48_clk),
    .Q(net54));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4799_ (.D(_0001_),
    .RN(net34),
    .CLK(clknet_leaf_48_clk),
    .Q(net55));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4800_ (.D(_0002_),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(net56));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4801_ (.D(_0003_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4802_ (.D(_0004_),
    .RN(net34),
    .CLK(clknet_leaf_48_clk),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4803_ (.D(_0005_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4804_ (.D(_0006_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4805_ (.D(_0007_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4806_ (.D(_0008_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4807_ (.D(_0009_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4808_ (.D(_0010_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4809_ (.D(_0011_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4810_ (.D(_0012_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4811_ (.D(_0013_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net70));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4812_ (.D(_0014_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net71));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4813_ (.D(_0015_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4814_ (.D(_0016_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net73));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4815_ (.D(_0017_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net74));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4816_ (.D(_0018_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net75));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4817_ (.D(_0019_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4818_ (.D(_0020_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4819_ (.D(_0021_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4820_ (.D(_0022_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4821_ (.D(_0023_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4822_ (.D(_0024_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4823_ (.D(_0025_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4824_ (.D(_0026_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4825_ (.D(_0027_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4826_ (.D(_0028_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[3].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4827_ (.D(_0029_),
    .RN(net34),
    .CLK(clknet_leaf_37_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4828_ (.D(_0030_),
    .RN(net34),
    .CLK(clknet_leaf_37_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4829_ (.D(_0031_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4830_ (.D(_0032_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4831_ (.D(_0033_),
    .RN(net34),
    .CLK(clknet_leaf_34_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4832_ (.D(_0034_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4833_ (.D(_0035_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4834_ (.D(_0036_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4835_ (.D(_0037_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4836_ (.D(_0038_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[13].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4837_ (.D(_0039_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4838_ (.D(_0040_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4839_ (.D(_0041_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4840_ (.D(_0042_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4841_ (.D(_0043_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4842_ (.D(_0044_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4843_ (.D(_0045_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4844_ (.D(_0046_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4845_ (.D(_0047_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4846_ (.D(_0048_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4847_ (.D(_0049_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4848_ (.D(_0050_),
    .RN(net34),
    .CLK(clknet_leaf_34_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4849_ (.D(_0051_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4850_ (.D(_0052_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4851_ (.D(_0053_),
    .RN(net34),
    .CLK(clknet_leaf_34_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4852_ (.D(_0054_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4853_ (.D(_0055_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4854_ (.D(_0056_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4855_ (.D(_0057_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4856_ (.D(\Stack_pointer.SP_next[0] ),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4857_ (.D(\Stack_pointer.SP_next[1] ),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4858_ (.D(\Stack_pointer.SP_next[2] ),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4859_ (.D(\Stack_pointer.SP_next[3] ),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(\Stack_pointer.SP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _4860_ (.D(\Stack_pointer.SP_next[4] ),
    .SETN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _4861_ (.D(\Stack_pointer.SP_next[5] ),
    .SETN(net34),
    .CLK(clknet_leaf_56_clk),
    .Q(\Stack_pointer.SP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _4862_ (.D(\Stack_pointer.SP_next[6] ),
    .SETN(net34),
    .CLK(clknet_leaf_56_clk),
    .Q(\Stack_pointer.SP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _4863_ (.D(\Stack_pointer.SP_next[7] ),
    .SETN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(\Stack_pointer.SP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4864_ (.D(_0058_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.p_Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4865_ (.D(\Control_unit1.instr_stage1[0] ),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_000.ALU_func[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4866_ (.D(\Control_unit1.instr_stage1[1] ),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_000.ALU_func[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4867_ (.D(\Control_unit1.instr_stage1[2] ),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4868_ (.D(\Control_unit1.instr_stage1[3] ),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(\Control_unit2.instr_stage2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4869_ (.D(\Control_unit1.instr_stage1[4] ),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(\Control_unit2.instr_stage2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4870_ (.D(\Control_unit1.instr_stage1[5] ),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(\Control_unit2.instr_stage2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4871_ (.D(\Control_unit1.instr_stage1[6] ),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(\Control_unit2.instr_stage2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4872_ (.D(\Control_unit1.instr_stage1[7] ),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(\Control_unit2.instr_stage2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4873_ (.D(\Control_unit1.instr_stage1[8] ),
    .RN(net34),
    .CLK(clknet_leaf_56_clk),
    .Q(\Control_unit2.instr_stage2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4874_ (.D(\Control_unit1.instr_stage1[9] ),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4875_ (.D(\Control_unit1.instr_stage1[10] ),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4876_ (.D(\Control_unit1.instr_stage1[11] ),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4877_ (.D(\Control_unit1.instr_stage1[12] ),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(\Control_unit2.instr_stage2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4878_ (.D(\Control_unit1.instr_decoder1.A[0] ),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(\Arithmetic_Logic_Unit.op ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _4879_ (.D(\Control_unit1.instr_decoder1.A[1] ),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4880_ (.D(\Control_unit1.instr_decoder1.A[2] ),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(\Control_unit2.instr_decoder2.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4881_ (.D(net2),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4882_ (.D(net9),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4883_ (.D(net10),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4884_ (.D(net11),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4885_ (.D(net12),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(\Control_unit1.instr_stage1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4886_ (.D(net13),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(\Control_unit1.instr_stage1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4887_ (.D(net14),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(\Control_unit1.instr_stage1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4888_ (.D(net15),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(\Control_unit1.instr_stage1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4889_ (.D(net16),
    .RN(net34),
    .CLK(clknet_leaf_56_clk),
    .Q(\Control_unit1.instr_stage1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4890_ (.D(net17),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(\Control_unit1.instr_stage1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4891_ (.D(net3),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(\Control_unit1.instr_stage1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4892_ (.D(net4),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(\Control_unit1.instr_stage1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4893_ (.D(net5),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(\Control_unit1.instr_stage1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4894_ (.D(net6),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4895_ (.D(net7),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(\Control_unit1.instr_decoder1.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4896_ (.D(net8),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(\Control_unit1.instr_decoder1.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4897_ (.D(_0059_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4898_ (.D(_0060_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4899_ (.D(_0061_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4900_ (.D(_0062_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4901_ (.D(_0063_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4902_ (.D(_0064_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4903_ (.D(_0065_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4904_ (.D(_0066_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4905_ (.D(_0067_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4906_ (.D(_0068_),
    .RN(net34),
    .CLK(clknet_leaf_34_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4907_ (.D(_0069_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4908_ (.D(_0070_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4909_ (.D(_0071_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4910_ (.D(_0072_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4911_ (.D(_0073_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4912_ (.D(_0074_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4913_ (.D(_0075_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4914_ (.D(_0076_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4915_ (.D(_0077_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4916_ (.D(_0078_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4917_ (.D(_0079_),
    .RN(net34),
    .CLK(clknet_leaf_43_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4918_ (.D(_0080_),
    .RN(net34),
    .CLK(clknet_leaf_43_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4919_ (.D(_0081_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4920_ (.D(_0082_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4921_ (.D(_0083_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4922_ (.D(_0084_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4923_ (.D(_0085_),
    .RN(net34),
    .CLK(clknet_leaf_26_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4924_ (.D(_0086_),
    .RN(net34),
    .CLK(clknet_leaf_26_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4925_ (.D(_0087_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4926_ (.D(_0088_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4927_ (.D(_0089_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4928_ (.D(_0090_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4929_ (.D(_0091_),
    .RN(net34),
    .CLK(clknet_leaf_62_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4930_ (.D(_0092_),
    .RN(net34),
    .CLK(clknet_leaf_62_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4931_ (.D(_0093_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4932_ (.D(_0094_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4933_ (.D(_0095_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4934_ (.D(_0096_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4935_ (.D(_0097_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4936_ (.D(_0098_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4937_ (.D(_0099_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4938_ (.D(_0100_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4939_ (.D(_0101_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4940_ (.D(_0102_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4941_ (.D(_0103_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4942_ (.D(_0104_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4943_ (.D(_0105_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4944_ (.D(_0106_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4945_ (.D(_0107_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4946_ (.D(_0108_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4947_ (.D(_0109_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4948_ (.D(_0110_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4949_ (.D(_0111_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4950_ (.D(_0112_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4951_ (.D(_0113_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4952_ (.D(_0114_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4953_ (.D(_0115_),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4954_ (.D(_0116_),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4955_ (.D(_0117_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4956_ (.D(_0118_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4957_ (.D(_0119_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4958_ (.D(_0120_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4959_ (.D(_0121_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4960_ (.D(_0122_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4961_ (.D(_0123_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4962_ (.D(_0124_),
    .RN(net34),
    .CLK(clknet_leaf_62_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4963_ (.D(_0125_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4964_ (.D(_0126_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4965_ (.D(_0127_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4966_ (.D(_0128_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4967_ (.D(_0129_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4968_ (.D(_0130_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4969_ (.D(_0131_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4970_ (.D(_0132_),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4971_ (.D(_0133_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4972_ (.D(_0134_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4973_ (.D(_0135_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4974_ (.D(_0136_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4975_ (.D(_0137_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4976_ (.D(_0138_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4977_ (.D(_0139_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4978_ (.D(_0140_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4979_ (.D(_0141_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4980_ (.D(_0142_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4981_ (.D(_0143_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4982_ (.D(_0144_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4983_ (.D(_0145_),
    .RN(net34),
    .CLK(clknet_leaf_14_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4984_ (.D(_0146_),
    .RN(net34),
    .CLK(clknet_leaf_14_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4985_ (.D(_0147_),
    .RN(net34),
    .CLK(clknet_leaf_20_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4986_ (.D(_0148_),
    .RN(net34),
    .CLK(clknet_leaf_20_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4987_ (.D(_0149_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4988_ (.D(_0150_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4989_ (.D(_0151_),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4990_ (.D(_0152_),
    .RN(net34),
    .CLK(clknet_leaf_7_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4991_ (.D(_0153_),
    .RN(net34),
    .CLK(clknet_leaf_7_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4992_ (.D(_0154_),
    .RN(net34),
    .CLK(clknet_leaf_7_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4993_ (.D(_0155_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4994_ (.D(_0156_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4995_ (.D(_0157_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4996_ (.D(_0158_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4997_ (.D(_0159_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4998_ (.D(_0160_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4999_ (.D(_0161_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5000_ (.D(_0162_),
    .RN(net34),
    .CLK(clknet_leaf_14_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5001_ (.D(_0163_),
    .RN(net34),
    .CLK(clknet_leaf_9_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5002_ (.D(_0164_),
    .RN(net34),
    .CLK(clknet_leaf_20_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5003_ (.D(_0165_),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5004_ (.D(_0166_),
    .RN(net34),
    .CLK(clknet_leaf_16_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5005_ (.D(_0167_),
    .RN(net34),
    .CLK(clknet_leaf_21_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5006_ (.D(_0168_),
    .RN(net34),
    .CLK(clknet_leaf_7_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5007_ (.D(_0169_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5008_ (.D(_0170_),
    .RN(net34),
    .CLK(clknet_leaf_7_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5009_ (.D(_0171_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5010_ (.D(_0172_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5011_ (.D(_0173_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5012_ (.D(_0174_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5013_ (.D(_0175_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5014_ (.D(_0176_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5015_ (.D(_0177_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5016_ (.D(_0178_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5017_ (.D(_0179_),
    .RN(net34),
    .CLK(clknet_leaf_9_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5018_ (.D(_0180_),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5019_ (.D(_0181_),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5020_ (.D(_0182_),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5021_ (.D(_0183_),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5022_ (.D(_0184_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5023_ (.D(_0185_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5024_ (.D(_0186_),
    .RN(net34),
    .CLK(clknet_leaf_7_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5025_ (.D(_0187_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5026_ (.D(_0188_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5027_ (.D(_0189_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5028_ (.D(_0190_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5029_ (.D(_0191_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5030_ (.D(_0192_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5031_ (.D(_0193_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5032_ (.D(_0194_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5033_ (.D(_0195_),
    .RN(net34),
    .CLK(clknet_leaf_9_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5034_ (.D(_0196_),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5035_ (.D(_0197_),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5036_ (.D(_0198_),
    .RN(net34),
    .CLK(clknet_leaf_9_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5037_ (.D(_0199_),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5038_ (.D(_0200_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5039_ (.D(_0201_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5040_ (.D(_0202_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5041_ (.D(_0203_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5042_ (.D(_0204_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5043_ (.D(_0205_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5044_ (.D(_0206_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5045_ (.D(_0207_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5046_ (.D(_0208_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5047_ (.D(_0209_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5048_ (.D(_0210_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5049_ (.D(_0211_),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5050_ (.D(_0212_),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5051_ (.D(_0213_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5052_ (.D(_0214_),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5053_ (.D(_0215_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5054_ (.D(_0216_),
    .RN(net34),
    .CLK(clknet_leaf_4_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5055_ (.D(_0217_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5056_ (.D(_0218_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5057_ (.D(_0219_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5058_ (.D(_0220_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5059_ (.D(_0221_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5060_ (.D(_0222_),
    .RN(net34),
    .CLK(clknet_leaf_88_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5061_ (.D(_0223_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5062_ (.D(_0224_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5063_ (.D(_0225_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5064_ (.D(_0226_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5065_ (.D(_0227_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5066_ (.D(_0228_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5067_ (.D(_0229_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5068_ (.D(_0230_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5069_ (.D(_0231_),
    .RN(net34),
    .CLK(clknet_leaf_2_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5070_ (.D(_0232_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5071_ (.D(_0233_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5072_ (.D(_0234_),
    .RN(net34),
    .CLK(clknet_leaf_5_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5073_ (.D(_0235_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5074_ (.D(_0236_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5075_ (.D(_0237_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5076_ (.D(_0238_),
    .RN(net34),
    .CLK(clknet_leaf_88_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5077_ (.D(_0239_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5078_ (.D(_0240_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5079_ (.D(_0241_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5080_ (.D(_0242_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5081_ (.D(_0243_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5082_ (.D(_0244_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5083_ (.D(_0245_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5084_ (.D(_0246_),
    .RN(net34),
    .CLK(clknet_leaf_2_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5085_ (.D(_0247_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5086_ (.D(_0248_),
    .RN(net34),
    .CLK(clknet_leaf_4_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5087_ (.D(_0249_),
    .RN(net34),
    .CLK(clknet_leaf_5_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5088_ (.D(_0250_),
    .RN(net34),
    .CLK(clknet_leaf_5_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5089_ (.D(_0251_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5090_ (.D(_0252_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5091_ (.D(_0253_),
    .RN(net34),
    .CLK(clknet_leaf_88_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5092_ (.D(_0254_),
    .RN(net34),
    .CLK(clknet_leaf_88_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5093_ (.D(_0255_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5094_ (.D(_0256_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5095_ (.D(_0257_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5096_ (.D(_0258_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5097_ (.D(_0259_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5098_ (.D(_0260_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5099_ (.D(_0261_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5100_ (.D(_0262_),
    .RN(net34),
    .CLK(clknet_leaf_2_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5101_ (.D(_0263_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5102_ (.D(_0264_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5103_ (.D(_0265_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5104_ (.D(_0266_),
    .RN(net34),
    .CLK(clknet_leaf_5_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5105_ (.D(_0267_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5106_ (.D(_0268_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5107_ (.D(_0269_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5108_ (.D(_0270_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5109_ (.D(_0271_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5110_ (.D(_0272_),
    .RN(net34),
    .CLK(clknet_leaf_99_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5111_ (.D(_0273_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5112_ (.D(_0274_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5113_ (.D(_0275_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5114_ (.D(_0276_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5115_ (.D(_0277_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5116_ (.D(_0278_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5117_ (.D(_0279_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5118_ (.D(_0280_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5119_ (.D(_0281_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5120_ (.D(_0282_),
    .RN(net34),
    .CLK(clknet_leaf_107_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5121_ (.D(_0283_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5122_ (.D(_0284_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5123_ (.D(_0285_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5124_ (.D(_0286_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5125_ (.D(_0287_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5126_ (.D(_0288_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5127_ (.D(_0289_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5128_ (.D(_0290_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5129_ (.D(_0291_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5130_ (.D(_0292_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5131_ (.D(_0293_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5132_ (.D(_0294_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5133_ (.D(_0295_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5134_ (.D(_0296_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5135_ (.D(_0297_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5136_ (.D(_0298_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5137_ (.D(_0299_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5138_ (.D(_0300_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5139_ (.D(_0301_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5140_ (.D(_0302_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5141_ (.D(_0303_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5142_ (.D(_0304_),
    .RN(net34),
    .CLK(clknet_leaf_99_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5143_ (.D(_0305_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5144_ (.D(_0306_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5145_ (.D(_0307_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5146_ (.D(_0308_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5147_ (.D(_0309_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5148_ (.D(_0310_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5149_ (.D(_0311_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5150_ (.D(_0312_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5151_ (.D(_0313_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5152_ (.D(_0314_),
    .RN(net34),
    .CLK(clknet_leaf_107_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5153_ (.D(_0315_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5154_ (.D(_0316_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5155_ (.D(_0317_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5156_ (.D(_0318_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5157_ (.D(_0319_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5158_ (.D(_0320_),
    .RN(net34),
    .CLK(clknet_leaf_99_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5159_ (.D(_0321_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5160_ (.D(_0322_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5161_ (.D(_0323_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5162_ (.D(_0324_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5163_ (.D(_0325_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5164_ (.D(_0326_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5165_ (.D(_0327_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5166_ (.D(_0328_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5167_ (.D(_0329_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5168_ (.D(_0330_),
    .RN(net34),
    .CLK(clknet_leaf_107_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5169_ (.D(_0331_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5170_ (.D(_0332_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5171_ (.D(_0333_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5172_ (.D(_0334_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5173_ (.D(_0335_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5174_ (.D(_0336_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5175_ (.D(_0337_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5176_ (.D(_0338_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5177_ (.D(_0339_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5178_ (.D(_0340_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5179_ (.D(_0341_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5180_ (.D(_0342_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5181_ (.D(_0343_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5182_ (.D(_0344_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5183_ (.D(_0345_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5184_ (.D(_0346_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5185_ (.D(_0347_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5186_ (.D(_0348_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5187_ (.D(_0349_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5188_ (.D(_0350_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5189_ (.D(_0351_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5190_ (.D(_0352_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5191_ (.D(_0353_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5192_ (.D(_0354_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5193_ (.D(_0355_),
    .RN(net34),
    .CLK(clknet_leaf_99_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5194_ (.D(_0356_),
    .RN(net34),
    .CLK(clknet_leaf_99_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5195_ (.D(_0357_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5196_ (.D(_0358_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5197_ (.D(_0359_),
    .RN(net34),
    .CLK(clknet_leaf_2_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5198_ (.D(_0360_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5199_ (.D(_0361_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5200_ (.D(_0362_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5201_ (.D(_0363_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5202_ (.D(_0364_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5203_ (.D(_0365_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5204_ (.D(_0366_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5205_ (.D(_0367_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5206_ (.D(_0368_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5207_ (.D(_0369_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5208_ (.D(_0370_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5209_ (.D(_0371_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5210_ (.D(_0372_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5211_ (.D(_0373_),
    .RN(net34),
    .CLK(clknet_leaf_95_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5212_ (.D(_0374_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5213_ (.D(_0375_),
    .RN(net34),
    .CLK(clknet_leaf_2_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5214_ (.D(_0376_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5215_ (.D(_0377_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5216_ (.D(_0378_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5217_ (.D(_0379_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5218_ (.D(_0380_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5219_ (.D(_0381_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5220_ (.D(_0382_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5221_ (.D(_0383_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5222_ (.D(_0384_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5223_ (.D(_0385_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5224_ (.D(_0386_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5225_ (.D(_0387_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5226_ (.D(_0388_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5227_ (.D(_0389_),
    .RN(net34),
    .CLK(clknet_leaf_95_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5228_ (.D(_0390_),
    .RN(net34),
    .CLK(clknet_leaf_95_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5229_ (.D(_0391_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5230_ (.D(_0392_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5231_ (.D(_0393_),
    .RN(net34),
    .CLK(clknet_leaf_107_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5232_ (.D(_0394_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5233_ (.D(_0395_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5234_ (.D(_0396_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5235_ (.D(_0397_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5236_ (.D(_0398_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5237_ (.D(_0399_),
    .RN(net34),
    .CLK(clknet_leaf_89_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5238_ (.D(_0400_),
    .RN(net34),
    .CLK(clknet_leaf_89_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5239_ (.D(_0401_),
    .RN(net34),
    .CLK(clknet_leaf_89_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5240_ (.D(_0402_),
    .RN(net34),
    .CLK(clknet_leaf_89_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5241_ (.D(_0403_),
    .RN(net34),
    .CLK(clknet_leaf_95_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5242_ (.D(_0404_),
    .RN(net34),
    .CLK(clknet_leaf_95_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5243_ (.D(_0405_),
    .RN(net34),
    .CLK(clknet_leaf_95_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5244_ (.D(_0406_),
    .RN(net34),
    .CLK(clknet_leaf_95_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5245_ (.D(_0407_),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5246_ (.D(_0408_),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5247_ (.D(_0409_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5248_ (.D(_0410_),
    .RN(net34),
    .CLK(clknet_leaf_4_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5249_ (.D(_0411_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5250_ (.D(_0412_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5251_ (.D(_0413_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5252_ (.D(_0414_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5253_ (.D(_0415_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5254_ (.D(_0416_),
    .RN(net34),
    .CLK(clknet_leaf_89_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5255_ (.D(_0417_),
    .RN(net34),
    .CLK(clknet_leaf_89_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5256_ (.D(_0418_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5257_ (.D(_0419_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5258_ (.D(_0420_),
    .RN(net34),
    .CLK(clknet_leaf_95_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5259_ (.D(_0421_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5260_ (.D(_0422_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5261_ (.D(_0423_),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5262_ (.D(_0424_),
    .RN(net34),
    .CLK(clknet_leaf_10_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5263_ (.D(_0425_),
    .RN(net34),
    .CLK(clknet_leaf_10_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5264_ (.D(_0426_),
    .RN(net34),
    .CLK(clknet_leaf_4_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5265_ (.D(_0427_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5266_ (.D(_0428_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5267_ (.D(_0429_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5268_ (.D(_0430_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5269_ (.D(_0431_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5270_ (.D(_0432_),
    .RN(net34),
    .CLK(clknet_leaf_89_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5271_ (.D(_0433_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5272_ (.D(_0434_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5273_ (.D(_0435_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5274_ (.D(_0436_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5275_ (.D(_0437_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5276_ (.D(_0438_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5277_ (.D(_0439_),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5278_ (.D(_0440_),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5279_ (.D(_0441_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5280_ (.D(_0442_),
    .RN(net34),
    .CLK(clknet_leaf_10_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5281_ (.D(_0443_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5282_ (.D(_0444_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5283_ (.D(_0445_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5284_ (.D(_0446_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5285_ (.D(_0447_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5286_ (.D(_0448_),
    .RN(net34),
    .CLK(clknet_leaf_89_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5287_ (.D(_0449_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5288_ (.D(_0450_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5289_ (.D(_0451_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5290_ (.D(_0452_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5291_ (.D(_0453_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5292_ (.D(_0454_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5293_ (.D(_0455_),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5294_ (.D(_0456_),
    .RN(net34),
    .CLK(clknet_leaf_10_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5295_ (.D(_0457_),
    .RN(net34),
    .CLK(clknet_leaf_10_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5296_ (.D(_0458_),
    .RN(net34),
    .CLK(clknet_leaf_10_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5297_ (.D(_0459_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5298_ (.D(_0460_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5299_ (.D(_0461_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5300_ (.D(_0462_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5301_ (.D(_0463_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5302_ (.D(_0464_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5303_ (.D(_0465_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5304_ (.D(_0466_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5305_ (.D(_0467_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5306_ (.D(_0468_),
    .RN(net34),
    .CLK(clknet_leaf_14_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5307_ (.D(_0469_),
    .RN(net34),
    .CLK(clknet_leaf_16_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5308_ (.D(_0470_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5309_ (.D(_0471_),
    .RN(net34),
    .CLK(clknet_leaf_21_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5310_ (.D(_0472_),
    .RN(net34),
    .CLK(clknet_leaf_21_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5311_ (.D(_0473_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5312_ (.D(_0474_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5313_ (.D(_0475_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5314_ (.D(_0476_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5315_ (.D(_0477_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5316_ (.D(_0478_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5317_ (.D(_0479_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5318_ (.D(_0480_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5319_ (.D(_0481_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5320_ (.D(_0482_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5321_ (.D(_0483_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5322_ (.D(_0484_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5323_ (.D(_0485_),
    .RN(net34),
    .CLK(clknet_leaf_16_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5324_ (.D(_0486_),
    .RN(net34),
    .CLK(clknet_leaf_16_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5325_ (.D(_0487_),
    .RN(net34),
    .CLK(clknet_leaf_20_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5326_ (.D(_0488_),
    .RN(net34),
    .CLK(clknet_leaf_21_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5327_ (.D(_0489_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5328_ (.D(_0490_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5329_ (.D(_0491_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5330_ (.D(_0492_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5331_ (.D(_0493_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5332_ (.D(_0494_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5333_ (.D(_0495_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5334_ (.D(_0496_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5335_ (.D(_0497_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5336_ (.D(_0498_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5337_ (.D(_0499_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5338_ (.D(_0500_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5339_ (.D(_0501_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5340_ (.D(_0502_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5341_ (.D(_0503_),
    .RN(net34),
    .CLK(clknet_leaf_21_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5342_ (.D(_0504_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5343_ (.D(_0505_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5344_ (.D(_0506_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5345_ (.D(_0507_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5346_ (.D(_0508_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5347_ (.D(_0509_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5348_ (.D(_0510_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5349_ (.D(_0511_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5350_ (.D(_0512_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5351_ (.D(_0513_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5352_ (.D(_0514_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5353_ (.D(_0515_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5354_ (.D(_0516_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5355_ (.D(_0517_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5356_ (.D(_0518_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5357_ (.D(_0519_),
    .RN(net34),
    .CLK(clknet_leaf_21_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5358_ (.D(_0520_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5359_ (.D(_0521_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5360_ (.D(_0522_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5361_ (.D(_0523_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5362_ (.D(_0524_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5363_ (.D(_0525_),
    .RN(net34),
    .CLK(clknet_leaf_62_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5364_ (.D(_0526_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5365_ (.D(_0527_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5366_ (.D(_0528_),
    .RN(net34),
    .CLK(clknet_leaf_44_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5367_ (.D(_0529_),
    .RN(net34),
    .CLK(clknet_leaf_44_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5368_ (.D(_0530_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5369_ (.D(_0531_),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5370_ (.D(_0532_),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5371_ (.D(_0533_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5372_ (.D(_0534_),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5373_ (.D(_0535_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5374_ (.D(_0536_),
    .RN(net34),
    .CLK(clknet_leaf_29_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5375_ (.D(_0537_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5376_ (.D(_0538_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5377_ (.D(_0539_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5378_ (.D(_0540_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5379_ (.D(_0541_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5380_ (.D(_0542_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5381_ (.D(_0543_),
    .RN(net34),
    .CLK(clknet_leaf_43_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5382_ (.D(_0544_),
    .RN(net34),
    .CLK(clknet_leaf_44_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5383_ (.D(_0545_),
    .RN(net34),
    .CLK(clknet_leaf_43_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5384_ (.D(_0546_),
    .RN(net34),
    .CLK(clknet_leaf_43_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5385_ (.D(_0547_),
    .RN(net34),
    .CLK(clknet_leaf_35_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5386_ (.D(_0548_),
    .RN(net34),
    .CLK(clknet_leaf_35_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5387_ (.D(_0549_),
    .RN(net34),
    .CLK(clknet_leaf_26_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5388_ (.D(_0550_),
    .RN(net34),
    .CLK(clknet_leaf_35_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5389_ (.D(_0551_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5390_ (.D(_0552_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5391_ (.D(_0553_),
    .RN(net34),
    .CLK(clknet_leaf_29_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5392_ (.D(_0554_),
    .RN(net34),
    .CLK(clknet_leaf_29_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5393_ (.D(_0555_),
    .RN(net34),
    .CLK(clknet_leaf_49_clk),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5394_ (.D(_0556_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5395_ (.D(_0557_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5396_ (.D(_0558_),
    .RN(net34),
    .CLK(clknet_leaf_49_clk),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(Serial_input),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(instr[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(instr[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(instr[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(instr[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(instr[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(instr[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(instr[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(instr[1]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(instr[2]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(instr[3]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(instr[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(instr[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(instr[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(instr[7]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(instr[8]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(instr[9]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(read_data[0]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(read_data[10]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(read_data[11]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input21 (.I(read_data[12]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input22 (.I(read_data[13]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(read_data[14]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(read_data[15]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input25 (.I(read_data[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input26 (.I(read_data[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input27 (.I(read_data[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(read_data[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(read_data[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input30 (.I(read_data[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input31 (.I(read_data[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input32 (.I(read_data[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input33 (.I(read_data[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input34 (.I(reset),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(start),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output36 (.I(net36),
    .Z(Dataw_en));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output37 (.I(net37),
    .Z(Serial_output));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output38 (.I(net38),
    .Z(data_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output39 (.I(net39),
    .Z(data_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output40 (.I(net40),
    .Z(data_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output41 (.I(net41),
    .Z(data_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output42 (.I(net42),
    .Z(data_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output43 (.I(net43),
    .Z(data_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output44 (.I(net44),
    .Z(data_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output45 (.I(net45),
    .Z(data_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output46 (.I(net46),
    .Z(hlt));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output47 (.I(net47),
    .Z(instr_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output48 (.I(net48),
    .Z(instr_mem_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output49 (.I(net49),
    .Z(instr_mem_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output50 (.I(net50),
    .Z(instr_mem_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output51 (.I(net51),
    .Z(instr_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output52 (.I(net52),
    .Z(instr_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output53 (.I(net53),
    .Z(instr_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output54 (.I(net54),
    .Z(instr_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output55 (.I(net55),
    .Z(instr_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output56 (.I(net56),
    .Z(instr_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output57 (.I(net57),
    .Z(instr_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output58 (.I(net58),
    .Z(instr_mem_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output59 (.I(net59),
    .Z(instr_mem_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output60 (.I(net60),
    .Z(write_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output61 (.I(net61),
    .Z(write_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output62 (.I(net62),
    .Z(write_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output63 (.I(net63),
    .Z(write_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output64 (.I(net64),
    .Z(write_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output65 (.I(net65),
    .Z(write_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output66 (.I(net66),
    .Z(write_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output67 (.I(net67),
    .Z(write_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output68 (.I(net68),
    .Z(write_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output69 (.I(net69),
    .Z(write_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output70 (.I(net70),
    .Z(write_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output71 (.I(net71),
    .Z(write_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output72 (.I(net72),
    .Z(write_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output73 (.I(net73),
    .Z(write_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output74 (.I(net74),
    .Z(write_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output75 (.I(net75),
    .Z(write_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_opt_1_0_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_opt_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__B2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__B1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__B (.I(\Arithmetic_Logic_Unit.ALU_001.p_Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__I (.I(\Arithmetic_Logic_Unit.ALU_001.p_Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.p_Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__I (.I(\Arithmetic_Logic_Unit.op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__A1 (.I(\Arithmetic_Logic_Unit.op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__D (.I(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A1 (.I(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A1 (.I(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__I (.I(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__D (.I(\Control_unit1.instr_decoder1.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__A1 (.I(\Control_unit1.instr_decoder1.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__I (.I(\Control_unit1.instr_decoder1.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__A1 (.I(\Control_unit1.instr_decoder1.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(\Control_unit1.instr_decoder1.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__D (.I(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__A1 (.I(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__B (.I(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A1 (.I(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__D (.I(\Control_unit1.instr_stage1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A1 (.I(\Control_unit1.instr_stage1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__D (.I(\Control_unit1.instr_stage1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A2 (.I(\Control_unit1.instr_stage1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A2 (.I(\Control_unit1.instr_stage1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__D (.I(\Control_unit1.instr_stage1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A1 (.I(\Control_unit1.instr_stage1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A1 (.I(\Control_unit1.instr_stage1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__D (.I(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__A1 (.I(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A1 (.I(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A2 (.I(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__D (.I(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__B2 (.I(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A2 (.I(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__D (.I(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A1 (.I(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A1 (.I(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__D (.I(\Control_unit1.instr_stage1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A1 (.I(\Control_unit1.instr_stage1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A1 (.I(\Control_unit1.instr_stage1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__D (.I(\Control_unit1.instr_stage1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A1 (.I(\Control_unit1.instr_stage1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__A1 (.I(\Control_unit1.instr_stage1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__D (.I(\Control_unit1.instr_stage1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__A1 (.I(\Control_unit1.instr_stage1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A1 (.I(\Control_unit1.instr_stage1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__D (.I(\Control_unit1.instr_stage1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A1 (.I(\Control_unit1.instr_stage1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__A2 (.I(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__C (.I(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__I (.I(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A2 (.I(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__B (.I(\Control_unit2.instr_decoder2.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A1 (.I(\Control_unit2.instr_decoder2.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I (.I(\Control_unit2.instr_decoder2.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__I (.I(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A3 (.I(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A2 (.I(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__I (.I(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__I (.I(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__I (.I(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A2 (.I(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A2 (.I(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__I (.I(\Control_unit2.instr_stage2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__I (.I(\Control_unit2.instr_stage2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(\Control_unit2.instr_stage2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__A1 (.I(\Control_unit2.instr_stage2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(\Control_unit2.instr_stage2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A1 (.I(\Control_unit2.instr_stage2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(\Control_unit2.instr_stage2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A1 (.I(\Control_unit2.instr_stage2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A1 (.I(\Control_unit2.instr_stage2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A1 (.I(\Control_unit2.instr_stage2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A1 (.I(\Control_unit2.instr_stage2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A1 (.I(\Control_unit2.instr_stage2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A1 (.I(\Control_unit2.instr_stage2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__I (.I(\Control_unit2.instr_stage2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__I (.I(\Control_unit2.instr_stage2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__I (.I(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A2 (.I(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A1 (.I(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__I (.I(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(Serial_input));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__I (.I(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A1 (.I(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A1 (.I(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__B2 (.I(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A1 (.I(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A1 (.I(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__A1 (.I(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__C2 (.I(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A1 (.I(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A1 (.I(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__A1 (.I(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__B2 (.I(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A1 (.I(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A1 (.I(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A1 (.I(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__B2 (.I(\Stack_pointer.SP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A1 (.I(\Stack_pointer.SP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A1 (.I(\Stack_pointer.SP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__B2 (.I(\Stack_pointer.SP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A1 (.I(\Stack_pointer.SP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A1 (.I(\Stack_pointer.SP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__D (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__D (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__D (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__D (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__D (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__D (.I(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__D (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__D (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__D (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__D (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__D (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__D (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__I1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__C2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__B1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__I0 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__I1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__C2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__B1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__B1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__I0 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__B2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__I1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__I1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__B (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__B2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A3 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__I (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__B (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__I (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__A2 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__B (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__B1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__B1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__C (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__I (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__I (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__B1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__B1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__B1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__B1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__B (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__B (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__B1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__S (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__B (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__B1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__B1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__B1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__B1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__B1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__B1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__B1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A3 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A3 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A3 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__I (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__I (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__I (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__I (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__I (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__I (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__I0 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__I (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__I (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__I0 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__I0 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__I0 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__I (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__I (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__I0 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__I (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__I (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__I (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__I (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__I0 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__I0 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__I0 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__I0 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__I0 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__I (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__I (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__S (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__I (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__I (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__I (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__S (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__S (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__S (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__S (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__S (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__S (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__B (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__B (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__B2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A3 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A3 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A4 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__A4 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__B1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__I (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__I (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__I (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__I (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__B (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__I (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__I (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__I (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__I (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__I (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__I (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__I (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__I (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__I (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__I (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3356__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__I (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__I (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__I (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__I (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__I (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__I (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A2 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A2 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A2 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A2 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__I (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__I (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A2 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A2 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A2 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__I (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__I (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__I (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__I (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__I (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__I (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__I (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__I (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A2 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A2 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__I (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__I (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__I (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__I (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__I (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__B (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__B (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__I (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__C (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__I (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A3 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__A2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A4 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__I (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A2 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A2 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__I (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__I (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__B2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__B2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__B (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__B (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A1 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__B (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__C2 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__I (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__I (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__I (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__S (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__S (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__B2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__C2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__B2 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__B (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A2 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A2 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__I (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__I (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A1 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__I (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__I (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__I (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__I (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__C2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__B2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__I (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__B1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__B1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__I (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__I (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__C1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__C1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__C1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__C1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__A1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__I1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__B (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__S (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__S (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__I (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__I (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__I (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__I (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__I (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__B2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__B2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__B (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__C (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__I (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__I (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A3 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__C2 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__B2 (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__B2 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A2 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__B2 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B2 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__I (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__I (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A3 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A2 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A2 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__I (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A4 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__B2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__B1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__I (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__I (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__I (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__I (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__I (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__I (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__I0 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__I1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__B2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__B1 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__B2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__B2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__C1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__C1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__B1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__C1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__I1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__I (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__I (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__I (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__I (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__C (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__I (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A2 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__I (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A2 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A1 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__S (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__S (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A3 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__I1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__B2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__A2 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A2 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A2 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A2 (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__C1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__C1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__A1 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__A1 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__A1 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__I (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__I (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__I1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__B2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__C2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__I1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__B2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__B2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A3 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3174__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__I (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__B (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__B (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__C2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__I1 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__B2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A1 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__I (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__I (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__I (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__I1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B2 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A2 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__B1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A1 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__A1 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__A1 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__I (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__I1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__A1 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__I1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__C2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__B2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A3 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__C (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__I1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__C2 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A2 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__C (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(instr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(instr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(instr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(instr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(instr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(instr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(instr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(instr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(instr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(instr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(instr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(instr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(instr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(instr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(instr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(instr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(read_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(read_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(read_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(read_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(read_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(read_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(read_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(read_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(read_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(read_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(read_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(read_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(read_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(read_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(read_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(read_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(reset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(start));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__D (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__SETN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__SETN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__SETN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__SETN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__B (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__I0 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A3 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A3 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A4 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__CLK (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__CLK (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__CLK (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__CLK (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__CLK (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__CLK (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__CLK (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__CLK (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__CLK (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__CLK (.I(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__CLK (.I(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__CLK (.I(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__CLK (.I(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__CLK (.I(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__CLK (.I(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__CLK (.I(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__CLK (.I(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__CLK (.I(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__CLK (.I(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__CLK (.I(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__CLK (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__CLK (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__CLK (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__CLK (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__CLK (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__CLK (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__CLK (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__CLK (.I(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__CLK (.I(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__CLK (.I(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__CLK (.I(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__CLK (.I(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__CLK (.I(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__CLK (.I(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__CLK (.I(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__CLK (.I(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__CLK (.I(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__CLK (.I(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__CLK (.I(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__CLK (.I(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__CLK (.I(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__CLK (.I(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__CLK (.I(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__CLK (.I(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__CLK (.I(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__CLK (.I(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__CLK (.I(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__CLK (.I(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_3_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_3_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_3_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_3_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_3_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_3_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_3_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_3_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_opt_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
endmodule

