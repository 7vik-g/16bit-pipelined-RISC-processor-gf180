// This is the unpowered netlist.
module user_proj_example (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire net35;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net36;
 wire net55;
 wire net56;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net37;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net57;
 wire net58;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net59;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net60;
 wire net61;
 wire \k.A[0][0] ;
 wire \k.A[0][1] ;
 wire \k.A[0][2] ;
 wire \k.A[0][3] ;
 wire \k.A[0][4] ;
 wire \k.A[0][5] ;
 wire \k.A[0][6] ;
 wire \k.A[0][7] ;
 wire \k.A[1][0] ;
 wire \k.A[1][1] ;
 wire \k.A[1][2] ;
 wire \k.A[1][3] ;
 wire \k.A[1][4] ;
 wire \k.A[1][5] ;
 wire \k.A[1][6] ;
 wire \k.A[1][7] ;
 wire \k.A[2][0] ;
 wire \k.A[2][1] ;
 wire \k.A[2][2] ;
 wire \k.A[2][3] ;
 wire \k.A[2][4] ;
 wire \k.A[2][5] ;
 wire \k.A[2][6] ;
 wire \k.A[2][7] ;
 wire \k.A[3][0] ;
 wire \k.A[3][1] ;
 wire \k.A[3][2] ;
 wire \k.A[3][3] ;
 wire \k.A[3][4] ;
 wire \k.A[3][5] ;
 wire \k.A[3][6] ;
 wire \k.A[3][7] ;
 wire \k.B[0][0] ;
 wire \k.B[0][1] ;
 wire \k.B[0][2] ;
 wire \k.B[0][3] ;
 wire \k.B[0][4] ;
 wire \k.B[0][5] ;
 wire \k.B[0][6] ;
 wire \k.B[0][7] ;
 wire \k.B[1][0] ;
 wire \k.B[1][1] ;
 wire \k.B[1][2] ;
 wire \k.B[1][3] ;
 wire \k.B[1][4] ;
 wire \k.B[1][5] ;
 wire \k.B[1][6] ;
 wire \k.B[1][7] ;
 wire \k.B[2][0] ;
 wire \k.B[2][1] ;
 wire \k.B[2][2] ;
 wire \k.B[2][3] ;
 wire \k.B[2][4] ;
 wire \k.B[2][5] ;
 wire \k.B[2][6] ;
 wire \k.B[2][7] ;
 wire \k.B[3][0] ;
 wire \k.B[3][1] ;
 wire \k.B[3][2] ;
 wire \k.B[3][3] ;
 wire \k.B[3][4] ;
 wire \k.B[3][5] ;
 wire \k.B[3][6] ;
 wire \k.B[3][7] ;
 wire net78;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net79;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net80;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net81;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net82;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net83;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net147;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net148;
 wire net176;
 wire net177;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3336_ (.I(\k.B[1][4] ),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3337_ (.A1(_0674_),
    .A2(\k.A[0][1] ),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3338_ (.I(\k.B[1][3] ),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3339_ (.I(_0696_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3340_ (.I(_0707_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3341_ (.I(\k.A[0][0] ),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3342_ (.A1(_0718_),
    .A2(_0729_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3343_ (.A1(_0685_),
    .A2(_0740_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3344_ (.I(\k.A[0][1] ),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3345_ (.A1(_0718_),
    .A2(_0762_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3346_ (.I(_0674_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3347_ (.I(_0784_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3348_ (.I(\k.A[0][0] ),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3349_ (.A1(_0795_),
    .A2(_0806_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3350_ (.A1(_0773_),
    .A2(_0817_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3351_ (.A1(_0828_),
    .A2(_0751_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3352_ (.I(\k.A[0][3] ),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3353_ (.I(\k.B[1][1] ),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3354_ (.I(_0861_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3355_ (.A1(_0850_),
    .A2(_0872_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3356_ (.I(\k.B[1][0] ),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3357_ (.I(_0894_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3358_ (.I(_0905_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3359_ (.I(\k.A[0][2] ),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3360_ (.I(_0927_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3361_ (.A1(_0916_),
    .A2(_0938_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3362_ (.I(\k.A[0][1] ),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3363_ (.I(\k.B[1][2] ),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3364_ (.I(_0971_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3365_ (.I(_0982_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3366_ (.A1(_0960_),
    .A2(_0993_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3367_ (.I(_0850_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3368_ (.I(_0872_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3369_ (.A1(_1015_),
    .A2(_0916_),
    .B1(_1026_),
    .B2(_0938_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3370_ (.A1(_0883_),
    .A2(_0949_),
    .B1(_1004_),
    .B2(_1037_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3371_ (.I(\k.A[0][4] ),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3372_ (.I(_1059_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3373_ (.I(\k.B[1][0] ),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3374_ (.A1(_1070_),
    .A2(_1081_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3375_ (.A1(_0927_),
    .A2(_0993_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3376_ (.A1(_1092_),
    .A2(_0883_),
    .A3(_1103_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3377_ (.A1(_1048_),
    .A2(_1114_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3378_ (.A1(_1048_),
    .A2(_1114_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3379_ (.A1(_0839_),
    .A2(_1125_),
    .B(_1136_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3380_ (.I(\k.B[1][5] ),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3381_ (.I(_1158_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3382_ (.A1(_1169_),
    .A2(_0729_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3383_ (.I(_0696_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3384_ (.A1(_1191_),
    .A2(\k.A[0][2] ),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3385_ (.A1(_1202_),
    .A2(_0685_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3386_ (.A1(_1180_),
    .A2(_1213_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3387_ (.I(\k.B[1][1] ),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3388_ (.A1(_1059_),
    .A2(_1235_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3389_ (.I(_0850_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3390_ (.I(_1081_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3391_ (.A1(_1257_),
    .A2(_1268_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3392_ (.I(_1070_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3393_ (.I(_1235_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3394_ (.A1(_1290_),
    .A2(_1268_),
    .B1(_1301_),
    .B2(_1257_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3395_ (.A1(_1246_),
    .A2(_1279_),
    .B1(_1103_),
    .B2(_1312_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3396_ (.A1(\k.A[0][3] ),
    .A2(_0982_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3397_ (.I(\k.A[0][5] ),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3398_ (.A1(_1345_),
    .A2(_0894_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3399_ (.A1(_1246_),
    .A2(_1334_),
    .A3(_1356_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3400_ (.A1(_1323_),
    .A2(_1367_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3401_ (.A1(_1224_),
    .A2(_1378_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3402_ (.A1(_1147_),
    .A2(_1389_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3403_ (.A1(_0751_),
    .A2(_1400_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3404_ (.A1(_0839_),
    .A2(_1125_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3405_ (.I(_0927_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3406_ (.A1(_1026_),
    .A2(_1433_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3407_ (.I(_0916_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3408_ (.I(_0960_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3409_ (.A1(_1455_),
    .A2(_1466_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3410_ (.I(_0993_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3411_ (.A1(_0806_),
    .A2(_1488_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3412_ (.I(_1301_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3413_ (.I(_0938_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3414_ (.I(_0905_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3415_ (.A1(_1466_),
    .A2(_1510_),
    .B1(_1521_),
    .B2(_1532_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3416_ (.A1(_1444_),
    .A2(_1477_),
    .B1(_1499_),
    .B2(_1543_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3417_ (.A1(_1279_),
    .A2(_1444_),
    .A3(_1004_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3418_ (.A1(_1554_),
    .A2(_1565_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3419_ (.A1(_1554_),
    .A2(_1565_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3420_ (.A1(_0740_),
    .A2(_1576_),
    .B(_1587_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3421_ (.A1(_1422_),
    .A2(_1598_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3422_ (.I(_1026_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3423_ (.A1(_1466_),
    .A2(_1619_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3424_ (.A1(_0949_),
    .A2(_1630_),
    .A3(_1499_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3425_ (.I(_0729_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3426_ (.I(_1652_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3427_ (.I(_1455_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3428_ (.A1(_1663_),
    .A2(_1674_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3429_ (.A1(_1630_),
    .A2(_1641_),
    .A3(_1685_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3430_ (.A1(_0740_),
    .A2(_1554_),
    .A3(_1565_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3431_ (.A1(_1696_),
    .A2(_1707_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3432_ (.A1(_1411_),
    .A2(_1609_),
    .A3(_1718_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3433_ (.A1(_1147_),
    .A2(_1389_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3434_ (.A1(_0751_),
    .A2(_1400_),
    .B(_1740_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3435_ (.A1(_1323_),
    .A2(_1367_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3436_ (.A1(_1224_),
    .A2(_1378_),
    .B(_1762_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3437_ (.A1(_1158_),
    .A2(\k.A[0][1] ),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3438_ (.A1(_0674_),
    .A2(\k.A[0][2] ),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3439_ (.A1(_0696_),
    .A2(\k.A[0][3] ),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3440_ (.A1(_1795_),
    .A2(_1806_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3441_ (.A1(_1784_),
    .A2(_1817_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3442_ (.A1(_1345_),
    .A2(\k.B[1][1] ),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3443_ (.I(_1345_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3444_ (.A1(_1850_),
    .A2(_0894_),
    .B1(_1235_),
    .B2(_1059_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3445_ (.A1(_1092_),
    .A2(_1839_),
    .B1(_1861_),
    .B2(_1334_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3446_ (.A1(\k.A[0][4] ),
    .A2(_0971_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3447_ (.A1(\k.A[0][6] ),
    .A2(\k.B[1][0] ),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3448_ (.A1(_1839_),
    .A2(_1883_),
    .A3(_1893_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3449_ (.A1(_1872_),
    .A2(_1904_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3450_ (.A1(_1828_),
    .A2(_1915_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3451_ (.A1(_1795_),
    .A2(_0773_),
    .B1(_1213_),
    .B2(_1180_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3452_ (.I(\k.B[1][6] ),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3453_ (.I(_1948_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3454_ (.A1(_1959_),
    .A2(_0806_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3455_ (.A1(_1937_),
    .A2(_1970_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3456_ (.A1(_1773_),
    .A2(_1926_),
    .A3(_1981_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3457_ (.A1(_1751_),
    .A2(_1992_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3458_ (.A1(_1422_),
    .A2(_1598_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3459_ (.A1(_2014_),
    .A2(_1411_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3460_ (.A1(_2003_),
    .A2(_2025_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3461_ (.A1(_2003_),
    .A2(_2025_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3462_ (.A1(_1729_),
    .A2(_2036_),
    .B(_2047_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3463_ (.A1(_1751_),
    .A2(_1992_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3464_ (.I(_1948_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3465_ (.I(_2080_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3466_ (.I(_1663_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3467_ (.A1(_2091_),
    .A2(_2102_),
    .A3(_1937_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3468_ (.A1(_1773_),
    .A2(_1926_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3469_ (.A1(_1773_),
    .A2(_1926_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3470_ (.A1(_1981_),
    .A2(_2123_),
    .B(_2134_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3471_ (.A1(\k.B[1][4] ),
    .A2(\k.A[0][3] ),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3472_ (.A1(_1202_),
    .A2(_2156_),
    .B1(_1817_),
    .B2(_1784_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3473_ (.A1(\k.B[1][6] ),
    .A2(_0960_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3474_ (.A1(_2167_),
    .A2(_2178_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3475_ (.A1(\k.B[1][7] ),
    .A2(_0729_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3476_ (.A1(_2189_),
    .A2(_2200_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3477_ (.A1(_1872_),
    .A2(_1904_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3478_ (.A1(_1828_),
    .A2(_1915_),
    .B(_2222_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3479_ (.A1(\k.B[1][5] ),
    .A2(\k.A[0][2] ),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3480_ (.A1(\k.B[1][3] ),
    .A2(_1059_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3481_ (.A1(_2156_),
    .A2(_2255_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3482_ (.A1(_2244_),
    .A2(_2265_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3483_ (.A1(\k.A[0][6] ),
    .A2(\k.B[1][1] ),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3484_ (.I(\k.A[0][6] ),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3485_ (.A1(_2298_),
    .A2(_0894_),
    .B1(_0861_),
    .B2(_1345_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3486_ (.A1(_1356_),
    .A2(_2287_),
    .B1(_2309_),
    .B2(_1883_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3487_ (.A1(\k.A[0][5] ),
    .A2(\k.B[1][2] ),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3488_ (.A1(\k.A[0][7] ),
    .A2(\k.B[1][0] ),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3489_ (.A1(_2287_),
    .A2(_2331_),
    .A3(_2342_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3490_ (.A1(_2320_),
    .A2(_2353_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3491_ (.A1(_2276_),
    .A2(_2363_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3492_ (.A1(_2233_),
    .A2(_2374_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3493_ (.A1(_2211_),
    .A2(_2385_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3494_ (.A1(_2145_),
    .A2(_2396_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3495_ (.A1(_2112_),
    .A2(_2407_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3496_ (.A1(_2069_),
    .A2(_2417_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3497_ (.A1(_2069_),
    .A2(_2417_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3498_ (.A1(_2058_),
    .A2(_2427_),
    .B(_2438_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3499_ (.A1(_2112_),
    .A2(_2407_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3500_ (.A1(_2145_),
    .A2(_2396_),
    .B(_2458_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3501_ (.I(_2080_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3502_ (.I(_2479_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3503_ (.I(_0762_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3504_ (.I(_2499_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3505_ (.I(_2509_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3506_ (.A1(_2489_),
    .A2(_2519_),
    .A3(_2167_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3507_ (.A1(_2189_),
    .A2(_2200_),
    .B(_2530_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3508_ (.A1(_2233_),
    .A2(_2374_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3509_ (.A1(_2211_),
    .A2(_2385_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3510_ (.A1(_2550_),
    .A2(_2560_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3511_ (.I(\k.B[1][7] ),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3512_ (.A1(_2577_),
    .A2(_2499_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3513_ (.I(_0674_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3514_ (.A1(_2592_),
    .A2(_1070_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3515_ (.A1(_1806_),
    .A2(_2599_),
    .B1(_2265_),
    .B2(_2244_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3516_ (.A1(_1948_),
    .A2(_1433_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3517_ (.A1(_2607_),
    .A2(_2615_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3518_ (.A1(_2585_),
    .A2(_2623_),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3519_ (.I(_2331_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3520_ (.A1(_2287_),
    .A2(_2342_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3521_ (.A1(_2637_),
    .A2(_2644_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3522_ (.A1(_2320_),
    .A2(_2651_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3523_ (.A1(_2276_),
    .A2(_2363_),
    .B(_2657_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3524_ (.I(\k.A[0][7] ),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3525_ (.A1(_2671_),
    .A2(_0861_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3526_ (.A1(_1893_),
    .A2(_2678_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3527_ (.A1(_2637_),
    .A2(_2644_),
    .B(_2685_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3528_ (.A1(_2298_),
    .A2(_0971_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3529_ (.A1(_2678_),
    .A2(_2688_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3530_ (.A1(_2687_),
    .A2(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3531_ (.A1(_0696_),
    .A2(_1850_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3532_ (.A1(_1169_),
    .A2(_0850_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3533_ (.A1(_2599_),
    .A2(_2691_),
    .A3(_2692_),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3534_ (.A1(_2690_),
    .A2(_2693_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3535_ (.A1(_2665_),
    .A2(_2694_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3536_ (.A1(_2630_),
    .A2(_2695_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3537_ (.A1(_2569_),
    .A2(_2696_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3538_ (.A1(_2540_),
    .A2(_2697_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3539_ (.A1(_2468_),
    .A2(_2698_),
    .Z(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3540_ (.A1(_2468_),
    .A2(_2698_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3541_ (.A1(_2448_),
    .A2(_2699_),
    .B(_2700_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3542_ (.A1(_2569_),
    .A2(_2696_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3543_ (.A1(_2540_),
    .A2(_2697_),
    .B(_2702_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3544_ (.I(_2489_),
    .Z(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3545_ (.I(_1433_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3546_ (.I(_2705_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3547_ (.A1(_2704_),
    .A2(_2706_),
    .A3(_2607_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3548_ (.I(\k.B[1][7] ),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3549_ (.I(_2708_),
    .Z(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3550_ (.I(_2519_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3551_ (.A1(_2709_),
    .A2(_2710_),
    .A3(_2623_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3552_ (.A1(_2707_),
    .A2(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3553_ (.A1(_2665_),
    .A2(_2694_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3554_ (.A1(_2630_),
    .A2(_2695_),
    .B(_2713_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3555_ (.A1(_2577_),
    .A2(_2705_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3556_ (.A1(_2592_),
    .A2(_1850_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3557_ (.A1(_2599_),
    .A2(_2691_),
    .Z(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3558_ (.A1(_2255_),
    .A2(_2716_),
    .B1(_2717_),
    .B2(_2692_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3559_ (.I(_1015_),
    .Z(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3560_ (.A1(_1948_),
    .A2(_2719_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3561_ (.A1(_2718_),
    .A2(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3562_ (.A1(_2715_),
    .A2(_2721_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3563_ (.A1(_2690_),
    .A2(_2693_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3564_ (.A1(_2687_),
    .A2(_2689_),
    .B(_2723_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3565_ (.A1(_1158_),
    .A2(_1070_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3566_ (.I(_2298_),
    .Z(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3567_ (.A1(_0707_),
    .A2(_2726_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3568_ (.A1(_2716_),
    .A2(_2725_),
    .A3(_2727_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3569_ (.I(_2671_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3570_ (.A1(_2729_),
    .A2(_1488_),
    .A3(_2287_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3571_ (.A1(_2728_),
    .A2(_2730_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3572_ (.A1(_2724_),
    .A2(_2731_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3573_ (.A1(_2722_),
    .A2(_2732_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3574_ (.A1(_2714_),
    .A2(_2733_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3575_ (.A1(_2712_),
    .A2(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3576_ (.A1(_2703_),
    .A2(_2735_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3577_ (.A1(_2701_),
    .A2(_2736_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3578_ (.I(\k.A[1][1] ),
    .Z(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3579_ (.I(_2738_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3580_ (.I(_2739_),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3581_ (.I(_2740_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3582_ (.I(\k.B[3][1] ),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3583_ (.I(_2742_),
    .Z(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3584_ (.A1(_2741_),
    .A2(_2743_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3585_ (.I(\k.A[1][0] ),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3586_ (.I(_2745_),
    .Z(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3587_ (.I(\k.B[3][2] ),
    .Z(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3588_ (.I(_2747_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3589_ (.I(_2748_),
    .Z(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3590_ (.A1(_2746_),
    .A2(_2749_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3591_ (.I(\k.B[3][0] ),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3592_ (.I(_2751_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3593_ (.I(\k.A[1][2] ),
    .Z(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3594_ (.I(_2753_),
    .Z(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3595_ (.I(_2754_),
    .Z(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3596_ (.A1(_2752_),
    .A2(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3597_ (.A1(_2750_),
    .A2(_2756_),
    .A3(_2744_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3598_ (.I(_2746_),
    .Z(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3599_ (.I(_2752_),
    .Z(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3600_ (.I(_2759_),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3601_ (.A1(_2758_),
    .A2(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3602_ (.A1(_2744_),
    .A2(_2757_),
    .A3(_2761_),
    .Z(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3603_ (.I(\k.B[3][3] ),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3604_ (.I(_2763_),
    .Z(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3605_ (.I(\k.A[1][0] ),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3606_ (.A1(_2764_),
    .A2(_2765_),
    .A3(_2739_),
    .A4(_2749_),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3607_ (.I(_2766_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3608_ (.I(\k.A[1][3] ),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3609_ (.I(_2768_),
    .Z(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3610_ (.I(_2769_),
    .Z(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3611_ (.I(_2770_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3612_ (.I(\k.B[3][0] ),
    .Z(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3613_ (.I(_2772_),
    .Z(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3614_ (.I(_2773_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3615_ (.I(\k.B[3][1] ),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3616_ (.I(_2775_),
    .Z(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3617_ (.I(_2776_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3618_ (.I(_2754_),
    .Z(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3619_ (.A1(_2771_),
    .A2(_2774_),
    .A3(_2777_),
    .A4(_2778_),
    .Z(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3620_ (.I(\k.B[3][3] ),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3621_ (.I(_2780_),
    .Z(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3622_ (.I(_2781_),
    .Z(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3623_ (.I(_2749_),
    .Z(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3624_ (.I(_2783_),
    .Z(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3625_ (.A1(_2782_),
    .A2(_2758_),
    .B1(_2741_),
    .B2(_2784_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3626_ (.I(_2743_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3627_ (.A1(_2771_),
    .A2(_2759_),
    .B1(_2786_),
    .B2(_2778_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3628_ (.A1(_2767_),
    .A2(_2779_),
    .A3(_2785_),
    .A4(_2787_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3629_ (.A1(_2767_),
    .A2(_2785_),
    .B1(_2787_),
    .B2(_2779_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3630_ (.I(_2740_),
    .Z(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3631_ (.I(_2743_),
    .Z(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3632_ (.I(_2778_),
    .Z(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3633_ (.I(_2774_),
    .Z(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3634_ (.A1(_2790_),
    .A2(_2791_),
    .B1(_2792_),
    .B2(_2793_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3635_ (.I(_2755_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3636_ (.A1(_2793_),
    .A2(_2790_),
    .A3(_2791_),
    .A4(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3637_ (.A1(_2750_),
    .A2(_2794_),
    .B(_2796_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3638_ (.A1(_2788_),
    .A2(_2789_),
    .B(_2797_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3639_ (.A1(_2788_),
    .A2(_2797_),
    .A3(_2789_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3640_ (.A1(_2762_),
    .A2(_2798_),
    .B(_2799_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3641_ (.I(_2738_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3642_ (.A1(_2781_),
    .A2(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3643_ (.I(\k.B[3][4] ),
    .Z(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3644_ (.I(_2803_),
    .Z(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3645_ (.A1(_2804_),
    .A2(_2765_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3646_ (.I(_2753_),
    .Z(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3647_ (.A1(_2806_),
    .A2(_2747_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3648_ (.A1(_2802_),
    .A2(_2805_),
    .A3(_2807_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3649_ (.I(\k.A[1][4] ),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3650_ (.I(_2809_),
    .Z(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3651_ (.I(_2810_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3652_ (.A1(_2811_),
    .A2(_2751_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3653_ (.A1(_2769_),
    .A2(_2775_),
    .Z(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3654_ (.A1(_2812_),
    .A2(_2813_),
    .A3(_2766_),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3655_ (.A1(_2808_),
    .A2(_2814_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3656_ (.I(_2779_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3657_ (.A1(_2816_),
    .A2(_2788_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3658_ (.A1(_2815_),
    .A2(_2817_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3659_ (.A1(_2815_),
    .A2(_2817_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3660_ (.A1(_2800_),
    .A2(_2818_),
    .B(_2819_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3661_ (.I(_2811_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3662_ (.I(_2821_),
    .Z(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3663_ (.A1(_2813_),
    .A2(_2767_),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3664_ (.A1(_2822_),
    .A2(_2793_),
    .A3(_2823_),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3665_ (.A1(_2813_),
    .A2(_2767_),
    .B(_2824_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3666_ (.I(\k.B[3][5] ),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3667_ (.I(_2826_),
    .Z(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3668_ (.A1(_2827_),
    .A2(_2746_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3669_ (.A1(_2780_),
    .A2(_2806_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3670_ (.I(\k.A[1][3] ),
    .Z(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3671_ (.A1(_2830_),
    .A2(_2747_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3672_ (.A1(_2803_),
    .A2(_2801_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3673_ (.A1(_2829_),
    .A2(_2831_),
    .A3(_2832_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3674_ (.A1(_2828_),
    .A2(_2833_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3675_ (.I(\k.A[1][5] ),
    .Z(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3676_ (.A1(_2835_),
    .A2(_2772_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3677_ (.I(\k.B[3][4] ),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3678_ (.A1(_2837_),
    .A2(_2745_),
    .B1(_2738_),
    .B2(_2763_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3679_ (.A1(_2803_),
    .A2(_2763_),
    .A3(_2745_),
    .A4(_2738_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3680_ (.A1(_2807_),
    .A2(_2838_),
    .B(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3681_ (.A1(_2821_),
    .A2(_2742_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3682_ (.A1(_2836_),
    .A2(_2840_),
    .A3(_2841_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3683_ (.A1(_2808_),
    .A2(_2814_),
    .Z(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3684_ (.A1(_2834_),
    .A2(_2842_),
    .A3(_2843_),
    .Z(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3685_ (.A1(_2825_),
    .A2(_2844_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3686_ (.A1(_2834_),
    .A2(_2842_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3687_ (.A1(_2834_),
    .A2(_2842_),
    .Z(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3688_ (.A1(_2846_),
    .A2(_2847_),
    .A3(_2843_),
    .B1(_2825_),
    .B2(_2844_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3689_ (.I(\k.B[3][6] ),
    .Z(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3690_ (.A1(_2849_),
    .A2(_2826_),
    .A3(\k.A[1][0] ),
    .A4(\k.A[1][1] ),
    .Z(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3691_ (.I(_2850_),
    .Z(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3692_ (.I(\k.B[3][6] ),
    .Z(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3693_ (.I(_2852_),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3694_ (.A1(_2853_),
    .A2(_2745_),
    .B1(_2801_),
    .B2(_2827_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3695_ (.A1(_2851_),
    .A2(_2854_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3696_ (.A1(_2809_),
    .A2(\k.B[3][2] ),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3697_ (.A1(\k.A[1][3] ),
    .A2(\k.B[3][3] ),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3698_ (.A1(_2837_),
    .A2(_2806_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3699_ (.A1(_2856_),
    .A2(_2857_),
    .A3(_2858_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3700_ (.A1(_2855_),
    .A2(_2859_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3701_ (.A1(_2828_),
    .A2(_2833_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3702_ (.I(\k.A[1][6] ),
    .Z(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3703_ (.I(_2862_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3704_ (.A1(_2863_),
    .A2(_2751_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3705_ (.A1(_2803_),
    .A2(_2801_),
    .B1(_2754_),
    .B2(_2763_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3706_ (.A1(_2858_),
    .A2(_2802_),
    .B1(_2865_),
    .B2(_2831_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3707_ (.I(_2835_),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3708_ (.A1(_2867_),
    .A2(_2776_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3709_ (.A1(_2864_),
    .A2(_2866_),
    .A3(_2868_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3710_ (.A1(_2860_),
    .A2(_2861_),
    .A3(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3711_ (.A1(_2840_),
    .A2(_2841_),
    .Z(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3712_ (.A1(_2840_),
    .A2(_2841_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3713_ (.A1(_2836_),
    .A2(_2871_),
    .B(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3714_ (.A1(_2846_),
    .A2(_2870_),
    .A3(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3715_ (.A1(_2848_),
    .A2(_2874_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3716_ (.A1(_2848_),
    .A2(_2874_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3717_ (.A1(_2820_),
    .A2(_2845_),
    .A3(_2875_),
    .B(_2876_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3718_ (.A1(_2840_),
    .A2(_2841_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3719_ (.A1(_2836_),
    .A2(_2871_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3720_ (.A1(_2878_),
    .A2(_2879_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3721_ (.A1(_2846_),
    .A2(_2870_),
    .Z(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3722_ (.A1(_2846_),
    .A2(_2870_),
    .Z(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3723_ (.A1(_2880_),
    .A2(_2881_),
    .B(_2882_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3724_ (.A1(_2860_),
    .A2(_2861_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3725_ (.A1(_2860_),
    .A2(_2861_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3726_ (.A1(_2869_),
    .A2(_2884_),
    .B(_2885_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3727_ (.A1(\k.A[1][3] ),
    .A2(\k.B[3][4] ),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3728_ (.A1(_2768_),
    .A2(_2780_),
    .B1(_2806_),
    .B2(_2837_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3729_ (.A1(_2829_),
    .A2(_2887_),
    .B1(_2888_),
    .B2(_2856_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3730_ (.A1(_2862_),
    .A2(_2775_),
    .Z(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3731_ (.A1(_2889_),
    .A2(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3732_ (.I(\k.A[1][7] ),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3733_ (.A1(_2892_),
    .A2(_2773_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3734_ (.A1(_2891_),
    .A2(_2893_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3735_ (.A1(_2851_),
    .A2(_2854_),
    .A3(_2859_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3736_ (.A1(\k.A[1][5] ),
    .A2(\k.B[3][2] ),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3737_ (.A1(\k.A[1][4] ),
    .A2(\k.B[3][3] ),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3738_ (.A1(_2887_),
    .A2(_2896_),
    .A3(_2897_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3739_ (.A1(_2849_),
    .A2(\k.A[1][1] ),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3740_ (.A1(\k.B[3][5] ),
    .A2(\k.A[1][2] ),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3741_ (.I(\k.B[3][7] ),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3742_ (.A1(_2901_),
    .A2(\k.A[1][0] ),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3743_ (.A1(_2899_),
    .A2(_2900_),
    .A3(_2902_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3744_ (.A1(_2850_),
    .A2(_2898_),
    .A3(_2903_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3745_ (.A1(_2895_),
    .A2(_2904_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3746_ (.A1(_2894_),
    .A2(_2905_),
    .Z(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3747_ (.A1(_2866_),
    .A2(_2868_),
    .Z(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3748_ (.A1(_2866_),
    .A2(_2868_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3749_ (.A1(_2864_),
    .A2(_2907_),
    .A3(_2908_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3750_ (.A1(_2907_),
    .A2(_2909_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3751_ (.A1(_2886_),
    .A2(_2906_),
    .A3(_2910_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3752_ (.A1(_2883_),
    .A2(_2911_),
    .Z(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3753_ (.A1(_2883_),
    .A2(_2911_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3754_ (.A1(_2877_),
    .A2(_2912_),
    .B(_2913_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3755_ (.A1(_2886_),
    .A2(_2906_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3756_ (.A1(_2886_),
    .A2(_2906_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3757_ (.A1(_2910_),
    .A2(_2915_),
    .B(_2916_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3758_ (.A1(_2889_),
    .A2(_2890_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3759_ (.A1(_2891_),
    .A2(_2893_),
    .B(_2918_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3760_ (.A1(_2895_),
    .A2(_2904_),
    .Z(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3761_ (.A1(_2894_),
    .A2(_2905_),
    .B(_2920_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3762_ (.I(_2837_),
    .Z(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3763_ (.A1(_2810_),
    .A2(_2922_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3764_ (.A1(_2887_),
    .A2(_2897_),
    .Z(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3765_ (.A1(_2857_),
    .A2(_2923_),
    .B1(_2924_),
    .B2(_2896_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3766_ (.I(_2892_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3767_ (.A1(_2926_),
    .A2(_2786_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3768_ (.A1(_2925_),
    .A2(_2927_),
    .Z(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3769_ (.I(_2898_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3770_ (.A1(_2851_),
    .A2(_2903_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3771_ (.A1(_2851_),
    .A2(_2903_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3772_ (.A1(_2929_),
    .A2(_2930_),
    .B(_2931_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3773_ (.A1(_2862_),
    .A2(_2748_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3774_ (.A1(_2867_),
    .A2(_2781_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3775_ (.A1(_2923_),
    .A2(_2933_),
    .A3(_2934_),
    .Z(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3776_ (.I(_2901_),
    .Z(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3777_ (.A1(_2936_),
    .A2(_2765_),
    .B1(_2739_),
    .B2(_2853_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3778_ (.A1(_2936_),
    .A2(_2853_),
    .A3(_2765_),
    .A4(_2739_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3779_ (.A1(_2900_),
    .A2(_2937_),
    .B(_2938_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3780_ (.A1(\k.B[3][7] ),
    .A2(\k.A[1][1] ),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3781_ (.A1(_2849_),
    .A2(_2753_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3782_ (.A1(_2768_),
    .A2(_2826_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3783_ (.A1(_2940_),
    .A2(_2941_),
    .A3(_2942_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3784_ (.A1(_2939_),
    .A2(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3785_ (.A1(_2935_),
    .A2(_2944_),
    .Z(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3786_ (.A1(_2932_),
    .A2(_2945_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3787_ (.A1(_2921_),
    .A2(_2928_),
    .A3(_2946_),
    .Z(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3788_ (.A1(_2919_),
    .A2(_2947_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3789_ (.A1(_2917_),
    .A2(_2948_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3790_ (.A1(_2917_),
    .A2(_2948_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3791_ (.A1(_2914_),
    .A2(_2949_),
    .B(_2950_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3792_ (.A1(_2928_),
    .A2(_2946_),
    .Z(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3793_ (.A1(_2921_),
    .A2(_2952_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3794_ (.A1(_2919_),
    .A2(_2947_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3795_ (.A1(_2953_),
    .A2(_2954_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3796_ (.I(_2926_),
    .Z(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3797_ (.I(_2956_),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3798_ (.I(_2777_),
    .Z(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3799_ (.I(_2958_),
    .Z(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3800_ (.A1(_2957_),
    .A2(_2959_),
    .A3(_2925_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3801_ (.A1(_2932_),
    .A2(_2945_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3802_ (.A1(_2928_),
    .A2(_2946_),
    .B(_2961_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3803_ (.A1(\k.A[1][5] ),
    .A2(\k.B[3][4] ),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3804_ (.A1(_2923_),
    .A2(_2934_),
    .Z(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3805_ (.A1(_2897_),
    .A2(_2963_),
    .B1(_2964_),
    .B2(_2933_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3806_ (.A1(_2939_),
    .A2(_2943_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3807_ (.A1(_2935_),
    .A2(_2944_),
    .B(_2966_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3808_ (.A1(\k.A[1][7] ),
    .A2(_2748_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3809_ (.A1(\k.A[1][6] ),
    .A2(_2780_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3810_ (.A1(_2963_),
    .A2(_2969_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3811_ (.A1(_2968_),
    .A2(_2970_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3812_ (.A1(\k.B[3][7] ),
    .A2(_2753_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3813_ (.A1(_2940_),
    .A2(_2941_),
    .Z(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3814_ (.A1(_2899_),
    .A2(_2972_),
    .B1(_2973_),
    .B2(_2942_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3815_ (.A1(_2809_),
    .A2(\k.B[3][5] ),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3816_ (.A1(_2830_),
    .A2(_2852_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3817_ (.A1(_2972_),
    .A2(_2975_),
    .A3(_2976_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3818_ (.A1(_2974_),
    .A2(_2977_),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3819_ (.A1(_2971_),
    .A2(_2978_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3820_ (.A1(_2967_),
    .A2(_2979_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3821_ (.A1(_2965_),
    .A2(_2980_),
    .Z(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3822_ (.A1(_2962_),
    .A2(_2981_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3823_ (.A1(_2960_),
    .A2(_2982_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3824_ (.A1(_2951_),
    .A2(_2955_),
    .A3(_2983_),
    .Z(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3825_ (.I(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3826_ (.A1(_2737_),
    .A2(_2985_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3827_ (.A1(_2917_),
    .A2(_2948_),
    .A3(_2914_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3828_ (.A1(_2468_),
    .A2(_2698_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3829_ (.A1(_2448_),
    .A2(_2988_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3830_ (.A1(_2987_),
    .A2(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3831_ (.A1(_2877_),
    .A2(_2912_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3832_ (.A1(_2877_),
    .A2(_2912_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3833_ (.A1(_2058_),
    .A2(_2427_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3834_ (.A1(_2820_),
    .A2(_2845_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3835_ (.A1(_1609_),
    .A2(_1718_),
    .B(_2014_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3836_ (.A1(_1411_),
    .A2(_2995_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3837_ (.A1(_2994_),
    .A2(_2996_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3838_ (.A1(_1685_),
    .A2(_2761_),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3839_ (.I(_2998_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3840_ (.I(_2746_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3841_ (.I(_3000_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3842_ (.I(_2790_),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3843_ (.A1(_3001_),
    .A2(_2760_),
    .A3(_3002_),
    .A4(_2958_),
    .Z(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3844_ (.I(_2760_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3845_ (.I(_3002_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3846_ (.A1(_3004_),
    .A2(_3005_),
    .B1(_2959_),
    .B2(_3001_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3847_ (.A1(_3003_),
    .A2(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3848_ (.I(_1510_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3849_ (.I(_3008_),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3850_ (.A1(_2102_),
    .A2(_3009_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3851_ (.I(_1674_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3852_ (.A1(_1663_),
    .A2(_3011_),
    .A3(_2509_),
    .A4(_3008_),
    .Z(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3853_ (.A1(_1477_),
    .A2(_3010_),
    .B(_3012_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3854_ (.A1(_3007_),
    .A2(_3013_),
    .Z(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3855_ (.A1(_3007_),
    .A2(_3013_),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3856_ (.A1(_2999_),
    .A2(_3014_),
    .B(_3015_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3857_ (.A1(_2757_),
    .A2(_3003_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3858_ (.A1(_1641_),
    .A2(_3012_),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3859_ (.A1(_3017_),
    .A2(_3018_),
    .Z(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3860_ (.A1(_3017_),
    .A2(_3018_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3861_ (.A1(_3016_),
    .A2(_3019_),
    .B(_3020_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3862_ (.A1(_2788_),
    .A2(_2789_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3863_ (.A1(_2797_),
    .A2(_3022_),
    .A3(_2762_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3864_ (.A1(_1696_),
    .A2(_1707_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3865_ (.A1(_3023_),
    .A2(_3024_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3866_ (.A1(_3023_),
    .A2(_3024_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3867_ (.A1(_3021_),
    .A2(_3025_),
    .B(_3026_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3868_ (.A1(_1422_),
    .A2(_1598_),
    .A3(_1718_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3869_ (.A1(_2815_),
    .A2(_2817_),
    .A3(_2800_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3870_ (.A1(_3028_),
    .A2(_3029_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3871_ (.A1(_3028_),
    .A2(_3029_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3872_ (.A1(_3027_),
    .A2(_3030_),
    .B(_3031_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3873_ (.A1(_1411_),
    .A2(_2994_),
    .A3(_2995_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3874_ (.A1(_3032_),
    .A2(_3033_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3875_ (.A1(_2997_),
    .A2(_3034_),
    .Z(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3876_ (.A1(_2820_),
    .A2(_2845_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3877_ (.A1(_2848_),
    .A2(_2874_),
    .A3(_3036_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3878_ (.I(_3037_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3879_ (.A1(_2003_),
    .A2(_2025_),
    .A3(_1729_),
    .Z(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3880_ (.A1(_3038_),
    .A2(_3039_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3881_ (.A1(_3038_),
    .A2(_3039_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3882_ (.A1(_3035_),
    .A2(_3040_),
    .B(_3041_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3883_ (.A1(_2991_),
    .A2(_2992_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3884_ (.A1(_2058_),
    .A2(_2427_),
    .A3(_3043_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3885_ (.A1(_2991_),
    .A2(_2992_),
    .A3(_2993_),
    .B1(_3042_),
    .B2(_3044_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3886_ (.A1(_2448_),
    .A2(_2988_),
    .A3(_2987_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3887_ (.A1(_3045_),
    .A2(_3046_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3888_ (.A1(_2701_),
    .A2(_2736_),
    .A3(_2985_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3889_ (.A1(_2990_),
    .A2(_3047_),
    .B(_3048_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3890_ (.A1(_2963_),
    .A2(_2969_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3891_ (.A1(_2968_),
    .A2(_2970_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3892_ (.A1(_3050_),
    .A2(_3051_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3893_ (.I(_2977_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3894_ (.A1(_2974_),
    .A2(_3053_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3895_ (.A1(_2971_),
    .A2(_2978_),
    .B(_3054_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3896_ (.A1(_2804_),
    .A2(_2863_),
    .B1(_2764_),
    .B2(\k.A[1][7] ),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3897_ (.A1(_2922_),
    .A2(\k.A[1][7] ),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3898_ (.A1(_2969_),
    .A2(_3057_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3899_ (.I(_3058_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3900_ (.A1(_3056_),
    .A2(_3059_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3901_ (.A1(_2936_),
    .A2(_2768_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3902_ (.A1(_2972_),
    .A2(_2976_),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3903_ (.A1(_2941_),
    .A2(_3061_),
    .B1(_3062_),
    .B2(_2975_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3904_ (.A1(_2826_),
    .A2(\k.A[1][5] ),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3905_ (.A1(\k.B[3][7] ),
    .A2(_2830_),
    .A3(_2849_),
    .A4(_2809_),
    .Z(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3906_ (.A1(_2901_),
    .A2(_2830_),
    .B1(_2852_),
    .B2(_2810_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3907_ (.A1(_3065_),
    .A2(_3066_),
    .Z(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3908_ (.A1(_3064_),
    .A2(_3067_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3909_ (.A1(_3063_),
    .A2(_3068_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3910_ (.A1(_3060_),
    .A2(_3069_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3911_ (.A1(_3055_),
    .A2(_3070_),
    .Z(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3912_ (.I(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3913_ (.A1(_3052_),
    .A2(_3072_),
    .Z(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3914_ (.A1(_2967_),
    .A2(_2979_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3915_ (.A1(_2965_),
    .A2(_2980_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3916_ (.A1(_3074_),
    .A2(_3075_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3917_ (.A1(_3073_),
    .A2(_3076_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3918_ (.A1(_2962_),
    .A2(_2981_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3919_ (.A1(_2960_),
    .A2(_2982_),
    .B(_3078_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3920_ (.A1(_3077_),
    .A2(_3079_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3921_ (.A1(_2953_),
    .A2(_2954_),
    .B(_2983_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3922_ (.A1(_2953_),
    .A2(_2954_),
    .A3(_2983_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3923_ (.A1(_2951_),
    .A2(_3081_),
    .B(_3082_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3924_ (.A1(_3080_),
    .A2(_3083_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3925_ (.A1(_2703_),
    .A2(_2735_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3926_ (.A1(_2701_),
    .A2(_2736_),
    .B(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3927_ (.A1(_2714_),
    .A2(_2733_),
    .Z(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3928_ (.A1(_2712_),
    .A2(_2734_),
    .B(_3087_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3929_ (.I(_2719_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3930_ (.I(_3089_),
    .Z(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3931_ (.A1(_2704_),
    .A2(_3090_),
    .A3(_2718_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3932_ (.I(_2706_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3933_ (.A1(_2709_),
    .A2(_3092_),
    .A3(_2721_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3934_ (.A1(_3091_),
    .A2(_3093_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3935_ (.A1(_2724_),
    .A2(_2731_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3936_ (.A1(_2722_),
    .A2(_2732_),
    .B(_3095_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3937_ (.A1(_2678_),
    .A2(_2688_),
    .B1(_2728_),
    .B2(_2730_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3938_ (.I(_1169_),
    .Z(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3939_ (.I(_1850_),
    .Z(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3940_ (.I(_3099_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3941_ (.A1(_3098_),
    .A2(_3100_),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3942_ (.A1(_0784_),
    .A2(_2726_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3943_ (.A1(_0707_),
    .A2(_2671_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3944_ (.A1(_3102_),
    .A2(_3103_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3945_ (.A1(_3101_),
    .A2(_3104_),
    .Z(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3946_ (.A1(_3097_),
    .A2(_3105_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3947_ (.A1(_2708_),
    .A2(_3089_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3948_ (.A1(_2716_),
    .A2(_2727_),
    .Z(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3949_ (.A1(_2691_),
    .A2(_3102_),
    .B1(_3108_),
    .B2(_2725_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3950_ (.I(_1290_),
    .Z(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3951_ (.A1(_1959_),
    .A2(_3110_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3952_ (.A1(_3109_),
    .A2(_3111_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3953_ (.A1(_3107_),
    .A2(_3112_),
    .Z(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3954_ (.A1(_3106_),
    .A2(_3113_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3955_ (.A1(_3096_),
    .A2(_3114_),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3956_ (.A1(_3094_),
    .A2(_3115_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3957_ (.A1(_3088_),
    .A2(_3116_),
    .Z(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3958_ (.A1(_3084_),
    .A2(_3086_),
    .A3(_3117_),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3959_ (.A1(_2986_),
    .A2(_3049_),
    .A3(_3118_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3960_ (.I(net16),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3961_ (.A1(net15),
    .A2(_3120_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3962_ (.I(_3121_),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3963_ (.I(_3122_),
    .Z(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3964_ (.A1(_2986_),
    .A2(_3049_),
    .B(_3118_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3965_ (.A1(_3119_),
    .A2(_3123_),
    .A3(_3124_),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3966_ (.I(\k.A[2][2] ),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3967_ (.A1(_2592_),
    .A2(_3126_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3968_ (.I(_0718_),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3969_ (.I(\k.A[2][1] ),
    .Z(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3970_ (.I(_3129_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3971_ (.A1(_3128_),
    .A2(_3130_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3972_ (.A1(_1191_),
    .A2(_3126_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3973_ (.A1(_0784_),
    .A2(\k.A[2][1] ),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3974_ (.A1(_3132_),
    .A2(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3975_ (.A1(_3098_),
    .A2(\k.A[2][0] ),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3976_ (.A1(_3127_),
    .A2(_3131_),
    .B1(_3134_),
    .B2(_3135_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3977_ (.I(\k.A[2][0] ),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3978_ (.I(_3137_),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3979_ (.A1(_2479_),
    .A2(_3138_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3980_ (.A1(_3136_),
    .A2(_3139_),
    .Z(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3981_ (.A1(_3135_),
    .A2(_3134_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3982_ (.I(\k.A[2][4] ),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3983_ (.A1(_3142_),
    .A2(_0872_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3984_ (.I(\k.A[2][3] ),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3985_ (.I(_3144_),
    .Z(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3986_ (.A1(_3145_),
    .A2(_1532_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3987_ (.I(\k.A[2][2] ),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3988_ (.A1(_3147_),
    .A2(_1488_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3989_ (.I(_3142_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3990_ (.I(\k.A[2][3] ),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3991_ (.A1(_3149_),
    .A2(_0916_),
    .B1(_1026_),
    .B2(_3150_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3992_ (.A1(_3143_),
    .A2(_3146_),
    .B1(_3148_),
    .B2(_3151_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3993_ (.A1(\k.A[2][3] ),
    .A2(_0982_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3994_ (.I(\k.A[2][5] ),
    .Z(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3995_ (.I(_3154_),
    .Z(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3996_ (.A1(_3155_),
    .A2(_0905_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3997_ (.A1(_3143_),
    .A2(_3153_),
    .A3(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3998_ (.A1(_3152_),
    .A2(_3157_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3999_ (.A1(_3152_),
    .A2(_3157_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4000_ (.A1(_3141_),
    .A2(_3158_),
    .B(_3159_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4001_ (.A1(_1169_),
    .A2(_3129_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4002_ (.I(\k.A[2][3] ),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4003_ (.A1(_3162_),
    .A2(_1191_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4004_ (.A1(_3127_),
    .A2(_3163_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4005_ (.A1(_3161_),
    .A2(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4006_ (.I(\k.A[2][4] ),
    .Z(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4007_ (.I(_3166_),
    .Z(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4008_ (.A1(_3167_),
    .A2(_1268_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4009_ (.I(_3154_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4010_ (.A1(_3169_),
    .A2(_1235_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4011_ (.I(_3142_),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4012_ (.A1(_3155_),
    .A2(_1268_),
    .B1(_1301_),
    .B2(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4013_ (.A1(_3168_),
    .A2(_3170_),
    .B1(_3172_),
    .B2(_3153_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4014_ (.A1(_3166_),
    .A2(_0982_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4015_ (.I(\k.A[2][6] ),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4016_ (.A1(_3175_),
    .A2(_0905_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4017_ (.A1(_3170_),
    .A2(_3174_),
    .A3(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4018_ (.A1(_3173_),
    .A2(_3177_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4019_ (.A1(_3165_),
    .A2(_3178_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4020_ (.A1(_3160_),
    .A2(_3179_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4021_ (.A1(_3160_),
    .A2(_3179_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4022_ (.A1(_3140_),
    .A2(_3180_),
    .B(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4023_ (.A1(_3162_),
    .A2(_2592_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4024_ (.A1(_3132_),
    .A2(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4025_ (.A1(_3161_),
    .A2(_3164_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4026_ (.A1(_3184_),
    .A2(_3185_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4027_ (.I(\k.A[2][1] ),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4028_ (.A1(_1959_),
    .A2(_3187_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4029_ (.I(\k.A[2][0] ),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4030_ (.A1(_2577_),
    .A2(_3189_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4031_ (.A1(_3186_),
    .A2(_3188_),
    .A3(_3190_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4032_ (.A1(_3173_),
    .A2(_3177_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4033_ (.A1(_3165_),
    .A2(_3178_),
    .B(_3192_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4034_ (.A1(_1158_),
    .A2(\k.A[2][2] ),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4035_ (.A1(_3171_),
    .A2(_1191_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4036_ (.A1(_3183_),
    .A2(_3194_),
    .A3(_3195_),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4037_ (.A1(\k.A[2][6] ),
    .A2(_0861_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4038_ (.A1(_3175_),
    .A2(_1081_),
    .B1(_0872_),
    .B2(_3169_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4039_ (.A1(_3156_),
    .A2(_3197_),
    .B1(_3198_),
    .B2(_3174_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4040_ (.A1(_3154_),
    .A2(_0971_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4041_ (.A1(\k.A[2][7] ),
    .A2(_1081_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4042_ (.A1(_3197_),
    .A2(_3200_),
    .A3(_3201_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4043_ (.A1(_3199_),
    .A2(_3202_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4044_ (.A1(_3196_),
    .A2(_3203_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4045_ (.A1(_3193_),
    .A2(_3204_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4046_ (.A1(_3191_),
    .A2(_3205_),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4047_ (.I(_3138_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4048_ (.I(_3207_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4049_ (.I(_3208_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4050_ (.A1(_2704_),
    .A2(_3209_),
    .A3(_3136_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4051_ (.A1(_3182_),
    .A2(_3206_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4052_ (.A1(_3210_),
    .A2(_3211_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4053_ (.A1(_3182_),
    .A2(_3206_),
    .B(_3212_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4054_ (.A1(_3186_),
    .A2(_3188_),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4055_ (.A1(_3186_),
    .A2(_3188_),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4056_ (.A1(_3214_),
    .A2(_3190_),
    .B(_3215_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4057_ (.A1(_3193_),
    .A2(_3204_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4058_ (.A1(_3191_),
    .A2(_3205_),
    .B(_3217_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4059_ (.A1(_3149_),
    .A2(_0795_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4060_ (.A1(_3183_),
    .A2(_3195_),
    .Z(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4061_ (.A1(_3163_),
    .A2(_3219_),
    .B1(_3220_),
    .B2(_3194_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4062_ (.I(_3147_),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4063_ (.A1(_1959_),
    .A2(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4064_ (.A1(_3221_),
    .A2(_3223_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4065_ (.I(_3130_),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4066_ (.A1(_2577_),
    .A2(_3225_),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4067_ (.A1(_3224_),
    .A2(_3226_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4068_ (.A1(_3199_),
    .A2(_3202_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4069_ (.A1(_3196_),
    .A2(_3203_),
    .B(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4070_ (.I(_3145_),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4071_ (.A1(_3230_),
    .A2(_3098_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4072_ (.I(_3155_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4073_ (.I(_3232_),
    .Z(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4074_ (.A1(_3233_),
    .A2(_3128_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4075_ (.A1(_3219_),
    .A2(_3231_),
    .A3(_3234_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4076_ (.I(\k.A[2][7] ),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4077_ (.I(_3236_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4078_ (.I(\k.A[2][6] ),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4079_ (.I(_3238_),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4080_ (.I(_3239_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4081_ (.A1(_3237_),
    .A2(_1455_),
    .B1(_1619_),
    .B2(_3240_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4082_ (.I(_3236_),
    .Z(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4083_ (.I(_3239_),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4084_ (.A1(_3242_),
    .A2(_3243_),
    .A3(_1455_),
    .A4(_1619_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4085_ (.A1(_3200_),
    .A2(_3241_),
    .B(_3244_),
    .ZN(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4086_ (.A1(_3242_),
    .A2(_1510_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4087_ (.I(_0993_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4088_ (.A1(_3243_),
    .A2(_3247_),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4089_ (.A1(_3246_),
    .A2(_3248_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4090_ (.A1(_3245_),
    .A2(_3249_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4091_ (.A1(_3235_),
    .A2(_3250_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4092_ (.A1(_3227_),
    .A2(_3229_),
    .A3(_3251_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4093_ (.A1(_3218_),
    .A2(_3252_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4094_ (.A1(_3216_),
    .A2(_3253_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4095_ (.A1(_0718_),
    .A2(_3137_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4096_ (.A1(_3133_),
    .A2(_3255_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4097_ (.I(_0795_),
    .Z(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4098_ (.A1(_3257_),
    .A2(_3189_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4099_ (.A1(_3131_),
    .A2(_3258_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4100_ (.A1(_3259_),
    .A2(_3256_),
    .ZN(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4101_ (.A1(_3144_),
    .A2(_1301_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4102_ (.A1(_1532_),
    .A2(_3222_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4103_ (.A1(_3187_),
    .A2(_1488_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4104_ (.I(_3126_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4105_ (.A1(_3145_),
    .A2(_1532_),
    .B1(_1510_),
    .B2(_3264_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4106_ (.A1(_3261_),
    .A2(_3262_),
    .B1(_3263_),
    .B2(_3265_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4107_ (.A1(_3168_),
    .A2(_3261_),
    .A3(_3148_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4108_ (.A1(_3266_),
    .A2(_3267_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4109_ (.A1(_3266_),
    .A2(_3267_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4110_ (.A1(_3260_),
    .A2(_3268_),
    .B(_3269_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4111_ (.A1(_3141_),
    .A2(_3158_),
    .Z(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4112_ (.A1(_3270_),
    .A2(_3271_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4113_ (.A1(_3256_),
    .A2(_3272_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4114_ (.A1(_3260_),
    .A2(_3268_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4115_ (.A1(_1619_),
    .A2(_3222_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4116_ (.I(_3187_),
    .Z(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4117_ (.A1(_1674_),
    .A2(_3276_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4118_ (.A1(_3189_),
    .A2(_3247_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4119_ (.I(_3264_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4120_ (.A1(_3130_),
    .A2(_3008_),
    .B1(_3279_),
    .B2(_1674_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4121_ (.A1(_3275_),
    .A2(_3277_),
    .B1(_3278_),
    .B2(_3280_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4122_ (.A1(_3146_),
    .A2(_3275_),
    .A3(_3263_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4123_ (.A1(_3281_),
    .A2(_3282_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4124_ (.A1(_3281_),
    .A2(_3282_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4125_ (.A1(_3255_),
    .A2(_3283_),
    .B(_3284_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4126_ (.A1(_3274_),
    .A2(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4127_ (.A1(_3276_),
    .A2(_3008_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4128_ (.A1(_3262_),
    .A2(_3287_),
    .A3(_3278_),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4129_ (.A1(_3207_),
    .A2(_3011_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4130_ (.A1(_3287_),
    .A2(_3288_),
    .A3(_3289_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4131_ (.A1(_3255_),
    .A2(_3281_),
    .A3(_3282_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4132_ (.A1(_3290_),
    .A2(_3291_),
    .ZN(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4133_ (.A1(_3273_),
    .A2(_3286_),
    .A3(_3292_),
    .Z(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4134_ (.A1(_3270_),
    .A2(_3271_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4135_ (.A1(_3256_),
    .A2(_3272_),
    .B(_3294_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4136_ (.A1(_3160_),
    .A2(_3179_),
    .A3(_3140_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4137_ (.A1(_3295_),
    .A2(_3296_),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4138_ (.A1(_3274_),
    .A2(_3285_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4139_ (.A1(_3298_),
    .A2(_3273_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4140_ (.A1(_3297_),
    .A2(_3299_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4141_ (.A1(_3297_),
    .A2(_3299_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4142_ (.A1(_3293_),
    .A2(_3300_),
    .B(_3301_),
    .ZN(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4143_ (.A1(_3295_),
    .A2(_3296_),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4144_ (.A1(_3210_),
    .A2(_3211_),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4145_ (.A1(_3303_),
    .A2(_3304_),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4146_ (.A1(_3303_),
    .A2(_3304_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4147_ (.A1(_3302_),
    .A2(_3305_),
    .B(_3306_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4148_ (.A1(_3213_),
    .A2(_3254_),
    .A3(_3307_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4149_ (.I(\k.A[3][2] ),
    .Z(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4150_ (.A1(_2922_),
    .A2(_3309_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4151_ (.I(_2782_),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4152_ (.I(\k.A[3][1] ),
    .Z(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4153_ (.I(_3312_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4154_ (.A1(_3311_),
    .A2(_3313_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4155_ (.I(\k.A[3][2] ),
    .Z(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4156_ (.A1(_2764_),
    .A2(_3315_),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4157_ (.A1(_2804_),
    .A2(\k.A[3][1] ),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4158_ (.A1(_3316_),
    .A2(_3317_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4159_ (.I(_2827_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4160_ (.A1(_3319_),
    .A2(\k.A[3][0] ),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4161_ (.A1(_3310_),
    .A2(_3314_),
    .B1(_3318_),
    .B2(_3320_),
    .ZN(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4162_ (.I(_2852_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4163_ (.I(_3322_),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4164_ (.I(\k.A[3][0] ),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4165_ (.I(_3324_),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4166_ (.A1(_3323_),
    .A2(_3325_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4167_ (.A1(_3321_),
    .A2(_3326_),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4168_ (.A1(_3320_),
    .A2(_3318_),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4169_ (.I(\k.A[3][4] ),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4170_ (.I(_3329_),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4171_ (.A1(_3330_),
    .A2(_2742_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4172_ (.I(\k.A[3][3] ),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4173_ (.I(_3332_),
    .Z(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4174_ (.I(_3333_),
    .Z(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4175_ (.A1(_2752_),
    .A2(_3334_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4176_ (.I(_3309_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4177_ (.A1(_0064_),
    .A2(_2783_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4178_ (.I(_3330_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4179_ (.I(_3332_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4180_ (.A1(_0066_),
    .A2(_2752_),
    .B1(_2743_),
    .B2(_0067_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4181_ (.A1(_3331_),
    .A2(_3335_),
    .B1(_0065_),
    .B2(_0068_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4182_ (.I(\k.A[3][3] ),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4183_ (.A1(_2749_),
    .A2(_0070_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4184_ (.I(\k.A[3][5] ),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4185_ (.I(_0072_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4186_ (.A1(_0073_),
    .A2(_2772_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4187_ (.A1(_3331_),
    .A2(_0071_),
    .A3(_0074_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4188_ (.A1(_0069_),
    .A2(_0075_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4189_ (.A1(_0069_),
    .A2(_0075_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4190_ (.A1(_3328_),
    .A2(_0076_),
    .B(_0077_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(_3319_),
    .A2(_3312_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4192_ (.A1(_2781_),
    .A2(_0070_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4193_ (.A1(_3310_),
    .A2(_0080_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4194_ (.A1(_0079_),
    .A2(_0081_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4195_ (.A1(_0066_),
    .A2(_2773_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4196_ (.I(_0072_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4197_ (.A1(_0084_),
    .A2(_2775_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4198_ (.I(_3329_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4199_ (.A1(_0073_),
    .A2(_2773_),
    .B1(_2776_),
    .B2(_0086_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4200_ (.A1(_0083_),
    .A2(_0085_),
    .B1(_0087_),
    .B2(_0071_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4201_ (.A1(_3329_),
    .A2(_2748_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4202_ (.I(\k.A[3][6] ),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4203_ (.I(_0090_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4204_ (.A1(_0091_),
    .A2(_2751_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4205_ (.A1(_0085_),
    .A2(_0089_),
    .A3(_0092_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4206_ (.A1(_0088_),
    .A2(_0093_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4207_ (.A1(_0082_),
    .A2(_0094_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4208_ (.A1(_0078_),
    .A2(_0095_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4209_ (.A1(_0078_),
    .A2(_0095_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4210_ (.A1(_3327_),
    .A2(_0096_),
    .B(_0097_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4211_ (.A1(_2922_),
    .A2(_3332_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4212_ (.A1(_3316_),
    .A2(_0099_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4213_ (.A1(_0079_),
    .A2(_0081_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4214_ (.A1(_0100_),
    .A2(_0101_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4215_ (.I(\k.A[3][1] ),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4216_ (.A1(_3322_),
    .A2(_0103_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4217_ (.I(_2901_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4218_ (.I(\k.A[3][0] ),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4219_ (.A1(_0105_),
    .A2(_0106_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4220_ (.A1(_0102_),
    .A2(_0104_),
    .A3(_0107_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4221_ (.A1(_0088_),
    .A2(_0093_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4222_ (.A1(_0082_),
    .A2(_0094_),
    .B(_0109_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4223_ (.A1(_2827_),
    .A2(_3309_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4224_ (.A1(_2764_),
    .A2(_0086_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4225_ (.A1(_0099_),
    .A2(_0111_),
    .A3(_0112_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4226_ (.A1(\k.A[3][6] ),
    .A2(\k.B[3][1] ),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4227_ (.A1(_0091_),
    .A2(_2772_),
    .B1(_2742_),
    .B2(_0073_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4228_ (.A1(_0074_),
    .A2(_0114_),
    .B1(_0115_),
    .B2(_0089_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4229_ (.A1(_0072_),
    .A2(_2747_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4230_ (.A1(\k.A[3][7] ),
    .A2(\k.B[3][0] ),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4231_ (.A1(_0114_),
    .A2(_0117_),
    .A3(_0118_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4232_ (.A1(_0116_),
    .A2(_0119_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4233_ (.A1(_0113_),
    .A2(_0120_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4234_ (.A1(_0110_),
    .A2(_0121_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4235_ (.A1(_0108_),
    .A2(_0122_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4236_ (.I(_3323_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4237_ (.I(_0124_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4238_ (.I(_3325_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4239_ (.I(_0126_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4240_ (.I(_0127_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4241_ (.A1(_0125_),
    .A2(_0128_),
    .A3(_3321_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4242_ (.A1(_0098_),
    .A2(_0123_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4243_ (.A1(_0129_),
    .A2(_0130_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4244_ (.A1(_0098_),
    .A2(_0123_),
    .B(_0131_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4245_ (.A1(_0102_),
    .A2(_0104_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4246_ (.A1(_0102_),
    .A2(_0104_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4247_ (.A1(_0133_),
    .A2(_0107_),
    .B(_0134_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4248_ (.A1(_0110_),
    .A2(_0121_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4249_ (.A1(_0108_),
    .A2(_0122_),
    .B(_0136_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4250_ (.I(_2804_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4251_ (.I(_0066_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4252_ (.A1(_0138_),
    .A2(_0139_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4253_ (.A1(_0099_),
    .A2(_0112_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4254_ (.A1(_0080_),
    .A2(_0140_),
    .B1(_0141_),
    .B2(_0111_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4255_ (.I(_0064_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4256_ (.A1(_3322_),
    .A2(_0143_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4257_ (.A1(_0142_),
    .A2(_0144_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4258_ (.I(_3313_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4259_ (.A1(_0105_),
    .A2(_0146_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4260_ (.A1(_0145_),
    .A2(_0147_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4261_ (.A1(_0116_),
    .A2(_0119_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4262_ (.A1(_0113_),
    .A2(_0120_),
    .B(_0149_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4263_ (.I(_3319_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4264_ (.A1(_0151_),
    .A2(_3334_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4265_ (.I(_0084_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4266_ (.I(_0153_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4267_ (.A1(_3311_),
    .A2(_0154_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4268_ (.A1(_0140_),
    .A2(_0152_),
    .A3(_0155_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4269_ (.I(\k.A[3][7] ),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4270_ (.I(_0157_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4271_ (.I(_0158_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4272_ (.I(_0090_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4273_ (.I(_0160_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4274_ (.I(_0161_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4275_ (.A1(_0159_),
    .A2(_2759_),
    .B1(_2786_),
    .B2(_0162_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4276_ (.A1(_0159_),
    .A2(_0162_),
    .A3(_2759_),
    .A4(_2786_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4277_ (.A1(_0117_),
    .A2(_0163_),
    .B(_0164_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4278_ (.A1(_0158_),
    .A2(_2777_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4279_ (.A1(_0161_),
    .A2(_2783_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4280_ (.A1(_0166_),
    .A2(_0167_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4281_ (.A1(_0165_),
    .A2(_0168_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4282_ (.A1(_0156_),
    .A2(_0169_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4283_ (.A1(_0148_),
    .A2(_0150_),
    .A3(_0170_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4284_ (.A1(_0137_),
    .A2(_0171_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4285_ (.A1(_0135_),
    .A2(_0172_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4286_ (.A1(_3311_),
    .A2(_0106_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4287_ (.A1(_3317_),
    .A2(_0174_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4288_ (.I(_0138_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4289_ (.A1(_0176_),
    .A2(_3325_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4290_ (.A1(_3314_),
    .A2(_0177_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4291_ (.A1(_0178_),
    .A2(_0175_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_2776_),
    .A2(_3333_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4293_ (.I(_3315_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4294_ (.A1(_2774_),
    .A2(_0181_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4295_ (.A1(_0103_),
    .A2(_2783_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4296_ (.A1(_2777_),
    .A2(_0181_),
    .B1(_3334_),
    .B2(_2774_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4297_ (.A1(_0180_),
    .A2(_0182_),
    .B1(_0183_),
    .B2(_0184_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4298_ (.A1(_0083_),
    .A2(_0180_),
    .A3(_0065_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4299_ (.A1(_0185_),
    .A2(_0186_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4300_ (.A1(_0185_),
    .A2(_0186_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4301_ (.A1(_0179_),
    .A2(_0187_),
    .B(_0188_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4302_ (.A1(_3328_),
    .A2(_0076_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4303_ (.A1(_0189_),
    .A2(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4304_ (.A1(_0175_),
    .A2(_0191_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4305_ (.A1(_0179_),
    .A2(_0187_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4306_ (.A1(_2791_),
    .A2(_0143_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4307_ (.I(_3313_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4308_ (.A1(_2760_),
    .A2(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4309_ (.A1(_0106_),
    .A2(_2784_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4310_ (.I(_0143_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4311_ (.A1(_3313_),
    .A2(_2791_),
    .B1(_0198_),
    .B2(_2793_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4312_ (.A1(_0194_),
    .A2(_0196_),
    .B1(_0197_),
    .B2(_0199_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4313_ (.A1(_3335_),
    .A2(_0194_),
    .A3(_0183_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4314_ (.A1(_0200_),
    .A2(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4315_ (.A1(_0200_),
    .A2(_0201_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4316_ (.A1(_0174_),
    .A2(_0202_),
    .B(_0203_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4317_ (.A1(_0193_),
    .A2(_0204_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4318_ (.A1(_0195_),
    .A2(_2958_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4319_ (.A1(_0182_),
    .A2(_0206_),
    .A3(_0197_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4320_ (.A1(_3004_),
    .A2(_0126_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4321_ (.A1(_0206_),
    .A2(_0207_),
    .A3(_0208_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4322_ (.A1(_0174_),
    .A2(_0200_),
    .A3(_0201_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4323_ (.A1(_0209_),
    .A2(_0210_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4324_ (.A1(_0205_),
    .A2(_0211_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4325_ (.A1(_0192_),
    .A2(_0212_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4326_ (.A1(_0189_),
    .A2(_0190_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4327_ (.A1(_0175_),
    .A2(_0191_),
    .B(_0214_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4328_ (.A1(_0078_),
    .A2(_0095_),
    .A3(_3327_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4329_ (.A1(_0215_),
    .A2(_0216_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4330_ (.A1(_0193_),
    .A2(_0204_),
    .A3(_0192_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4331_ (.A1(_0217_),
    .A2(_0218_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4332_ (.A1(_0217_),
    .A2(_0218_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4333_ (.A1(_0213_),
    .A2(_0219_),
    .B(_0220_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4334_ (.A1(_0215_),
    .A2(_0216_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4335_ (.A1(_0129_),
    .A2(_0130_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4336_ (.A1(_0222_),
    .A2(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4337_ (.A1(_0222_),
    .A2(_0223_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4338_ (.A1(_0221_),
    .A2(_0224_),
    .B(_0225_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4339_ (.A1(_0132_),
    .A2(_0173_),
    .A3(_0226_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4340_ (.A1(_3308_),
    .A2(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4341_ (.A1(_3302_),
    .A2(_3305_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4342_ (.A1(_0221_),
    .A2(_0224_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4343_ (.A1(_0229_),
    .A2(_0230_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4344_ (.A1(_3293_),
    .A2(_3300_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4345_ (.A1(_0213_),
    .A2(_0219_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4346_ (.A1(_3293_),
    .A2(_3300_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4347_ (.A1(_0213_),
    .A2(_0219_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4348_ (.A1(_0232_),
    .A2(_0233_),
    .A3(_0234_),
    .A4(_0235_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4349_ (.A1(_0232_),
    .A2(_0234_),
    .B1(_0235_),
    .B2(_0233_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4350_ (.A1(_3286_),
    .A2(_3292_),
    .B(_3298_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4351_ (.A1(_3273_),
    .A2(_0238_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4352_ (.A1(_0193_),
    .A2(_0204_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4353_ (.A1(_0205_),
    .A2(_0211_),
    .B(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4354_ (.A1(_0192_),
    .A2(_0241_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4355_ (.A1(_0239_),
    .A2(_0242_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4356_ (.A1(_3274_),
    .A2(_3285_),
    .A3(_3292_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4357_ (.A1(_0193_),
    .A2(_0204_),
    .A3(_0211_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4358_ (.A1(_0244_),
    .A2(_0245_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4359_ (.A1(_3290_),
    .A2(_3291_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4360_ (.A1(_0209_),
    .A2(_0210_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4361_ (.A1(_0247_),
    .A2(_0248_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4362_ (.A1(_3289_),
    .A2(_0208_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4363_ (.A1(_3208_),
    .A2(_3009_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4364_ (.I(_3225_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4365_ (.A1(_3207_),
    .A2(_3011_),
    .A3(_0252_),
    .A4(_3009_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4366_ (.A1(_3277_),
    .A2(_0251_),
    .B(_0253_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4367_ (.A1(_0126_),
    .A2(_2959_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4368_ (.I(_0146_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4369_ (.A1(_3004_),
    .A2(_0126_),
    .A3(_0256_),
    .A4(_2958_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4370_ (.A1(_0196_),
    .A2(_0255_),
    .B(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4371_ (.A1(_0254_),
    .A2(_0258_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4372_ (.A1(_0254_),
    .A2(_0258_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4373_ (.A1(_0250_),
    .A2(_0259_),
    .B(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4374_ (.A1(_3288_),
    .A2(_0253_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4375_ (.A1(_0207_),
    .A2(_0257_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4376_ (.A1(_0262_),
    .A2(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4377_ (.A1(_0262_),
    .A2(_0263_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4378_ (.A1(_0261_),
    .A2(_0264_),
    .B(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4379_ (.A1(_0247_),
    .A2(_0248_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4380_ (.A1(_0266_),
    .A2(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4381_ (.A1(_0244_),
    .A2(_0245_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4382_ (.A1(_0249_),
    .A2(_0268_),
    .B(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4383_ (.A1(_0246_),
    .A2(_0270_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4384_ (.A1(_0239_),
    .A2(_0242_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4385_ (.A1(_0271_),
    .A2(_0272_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4386_ (.A1(_0243_),
    .A2(_0273_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4387_ (.A1(_0237_),
    .A2(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4388_ (.A1(_0229_),
    .A2(_0230_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4389_ (.A1(_0231_),
    .A2(_0236_),
    .A3(_0275_),
    .B(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4390_ (.A1(_3308_),
    .A2(_0227_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4391_ (.A1(_0228_),
    .A2(_0277_),
    .B(_0278_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4392_ (.A1(_3213_),
    .A2(_3254_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4393_ (.A1(_3213_),
    .A2(_3254_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4394_ (.A1(_3307_),
    .A2(_0280_),
    .B(_0281_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4395_ (.A1(_3218_),
    .A2(_3252_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4396_ (.A1(_3216_),
    .A2(_3253_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4397_ (.I(_2489_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4398_ (.I(_3279_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4399_ (.A1(_0285_),
    .A2(_0286_),
    .A3(_3221_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4400_ (.A1(_3224_),
    .A2(_3226_),
    .B(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4401_ (.A1(_3229_),
    .A2(_3251_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4402_ (.A1(_3229_),
    .A2(_3251_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4403_ (.A1(_3227_),
    .A2(_0289_),
    .B(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4404_ (.I(_2708_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4405_ (.A1(_0292_),
    .A2(_0286_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4406_ (.A1(_3232_),
    .A2(_0784_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4407_ (.A1(_3219_),
    .A2(_3234_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4408_ (.A1(_3195_),
    .A2(_0294_),
    .B1(_0295_),
    .B2(_3231_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4409_ (.A1(_3230_),
    .A2(_2479_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4410_ (.A1(_0296_),
    .A2(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4411_ (.A1(_0293_),
    .A2(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4412_ (.A1(_3245_),
    .A2(_3249_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4413_ (.A1(_3235_),
    .A2(_3250_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4414_ (.A1(_0300_),
    .A2(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4415_ (.I(_3237_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4416_ (.A1(_0303_),
    .A2(_3247_),
    .A3(_3197_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4417_ (.I(_3098_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4418_ (.A1(_3149_),
    .A2(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4419_ (.A1(_3239_),
    .A2(_0707_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4420_ (.A1(_0294_),
    .A2(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4421_ (.A1(_0306_),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4422_ (.A1(_0304_),
    .A2(_0309_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4423_ (.A1(_0302_),
    .A2(_0310_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4424_ (.A1(_0299_),
    .A2(_0311_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4425_ (.A1(_0288_),
    .A2(_0291_),
    .A3(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4426_ (.A1(_0283_),
    .A2(_0284_),
    .B(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4427_ (.A1(_0283_),
    .A2(_0284_),
    .A3(_0313_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4428_ (.A1(_0314_),
    .A2(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4429_ (.A1(_0282_),
    .A2(_0316_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4430_ (.A1(_0132_),
    .A2(_0173_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4431_ (.A1(_0132_),
    .A2(_0173_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4432_ (.A1(_0226_),
    .A2(_0318_),
    .B(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4433_ (.A1(_0137_),
    .A2(_0171_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4434_ (.A1(_0135_),
    .A2(_0172_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4435_ (.I(_0198_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4436_ (.A1(_0125_),
    .A2(_0323_),
    .A3(_0142_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4437_ (.A1(_0145_),
    .A2(_0147_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4438_ (.A1(_0150_),
    .A2(_0170_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4439_ (.A1(_0150_),
    .A2(_0170_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4440_ (.A1(_0148_),
    .A2(_0326_),
    .B(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4441_ (.I(_0105_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4442_ (.A1(_0329_),
    .A2(_0198_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4443_ (.A1(_0138_),
    .A2(_0153_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4444_ (.A1(_0140_),
    .A2(_0155_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4445_ (.A1(_0112_),
    .A2(_0331_),
    .B1(_0332_),
    .B2(_0152_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4446_ (.I(_3334_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4447_ (.A1(_3323_),
    .A2(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4448_ (.A1(_0333_),
    .A2(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4449_ (.A1(_0330_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4450_ (.A1(_0165_),
    .A2(_0168_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4451_ (.A1(_0156_),
    .A2(_0169_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4452_ (.A1(_0338_),
    .A2(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4453_ (.I(_0159_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4454_ (.A1(_0341_),
    .A2(_2784_),
    .A3(_0114_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4455_ (.A1(_0151_),
    .A2(_0139_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4456_ (.A1(_2782_),
    .A2(_0160_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4457_ (.A1(_0331_),
    .A2(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4458_ (.A1(_0343_),
    .A2(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4459_ (.A1(_0342_),
    .A2(_0346_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4460_ (.A1(_0340_),
    .A2(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4461_ (.A1(_0337_),
    .A2(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4462_ (.A1(_0325_),
    .A2(_0328_),
    .A3(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4463_ (.A1(_0321_),
    .A2(_0322_),
    .B(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4464_ (.A1(_0321_),
    .A2(_0322_),
    .A3(_0350_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4465_ (.A1(_0351_),
    .A2(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4466_ (.A1(_0320_),
    .A2(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4467_ (.A1(_0317_),
    .A2(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4468_ (.A1(_0317_),
    .A2(_0354_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4469_ (.A1(_0279_),
    .A2(_0355_),
    .B(_0356_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4470_ (.A1(_0328_),
    .A2(_0349_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4471_ (.A1(_0328_),
    .A2(_0349_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4472_ (.A1(_0325_),
    .A2(_0358_),
    .B(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4473_ (.I(_0125_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4474_ (.I(_0334_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4475_ (.I(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4476_ (.A1(_0361_),
    .A2(_0363_),
    .A3(_0333_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4477_ (.I(_0329_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4478_ (.I(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4479_ (.A1(_0366_),
    .A2(_0323_),
    .A3(_0336_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4480_ (.A1(_0364_),
    .A2(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4481_ (.A1(_0340_),
    .A2(_0347_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4482_ (.A1(_0337_),
    .A2(_0348_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4483_ (.A1(_0369_),
    .A2(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4484_ (.A1(_0329_),
    .A2(_0362_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4485_ (.A1(_0138_),
    .A2(_0161_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4486_ (.A1(_0155_),
    .A2(_0373_),
    .B1(_0345_),
    .B2(_0343_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4487_ (.I(_0139_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4488_ (.A1(_3323_),
    .A2(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4489_ (.A1(_0374_),
    .A2(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4490_ (.A1(_0372_),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4491_ (.A1(_0166_),
    .A2(_0167_),
    .B1(_0342_),
    .B2(_0346_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4492_ (.A1(_0151_),
    .A2(_0154_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4493_ (.A1(_2782_),
    .A2(_0158_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4494_ (.A1(_0373_),
    .A2(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4495_ (.A1(_0380_),
    .A2(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4496_ (.A1(_0379_),
    .A2(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4497_ (.I(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4498_ (.A1(_0378_),
    .A2(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4499_ (.A1(_0371_),
    .A2(_0386_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4500_ (.A1(_0368_),
    .A2(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4501_ (.A1(_0360_),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4502_ (.A1(_0226_),
    .A2(_0318_),
    .B(_0351_),
    .C(_0319_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4503_ (.A1(_0352_),
    .A2(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4504_ (.A1(_0389_),
    .A2(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4505_ (.I(_0315_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4506_ (.A1(_0291_),
    .A2(_0312_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4507_ (.A1(_0291_),
    .A2(_0312_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4508_ (.A1(_0288_),
    .A2(_0394_),
    .B(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4509_ (.I(_3230_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4510_ (.I(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4511_ (.I(_0285_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4512_ (.A1(_0398_),
    .A2(_0399_),
    .A3(_0296_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4513_ (.I(_2709_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4514_ (.I(_0401_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4515_ (.I(_0286_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4516_ (.A1(_0402_),
    .A2(_0403_),
    .A3(_0298_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4517_ (.A1(_0400_),
    .A2(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4518_ (.A1(_0302_),
    .A2(_0310_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4519_ (.A1(_0299_),
    .A2(_0311_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4520_ (.A1(_0406_),
    .A2(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4521_ (.A1(_0397_),
    .A2(_0292_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4522_ (.A1(_3243_),
    .A2(_0795_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4523_ (.A1(_3234_),
    .A2(_0410_),
    .B1(_0308_),
    .B2(_0306_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4524_ (.I(_3149_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4525_ (.A1(_0412_),
    .A2(_2080_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4526_ (.A1(_0411_),
    .A2(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4527_ (.A1(_0409_),
    .A2(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4528_ (.A1(_3246_),
    .A2(_3248_),
    .B1(_0304_),
    .B2(_0309_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4529_ (.A1(_3233_),
    .A2(_0305_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4530_ (.A1(_3242_),
    .A2(_3128_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4531_ (.A1(_0410_),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4532_ (.A1(_0417_),
    .A2(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4533_ (.A1(_0416_),
    .A2(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4534_ (.A1(_0415_),
    .A2(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4535_ (.A1(_0408_),
    .A2(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4536_ (.A1(_0405_),
    .A2(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4537_ (.A1(_0396_),
    .A2(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4538_ (.I(_0314_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4539_ (.A1(_3307_),
    .A2(_0280_),
    .B(_0426_),
    .C(_0281_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4540_ (.A1(_0393_),
    .A2(_0425_),
    .A3(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4541_ (.A1(_0393_),
    .A2(_0427_),
    .B(_0425_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4542_ (.A1(_0428_),
    .A2(_0429_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4543_ (.A1(_0392_),
    .A2(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4544_ (.A1(_0357_),
    .A2(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4545_ (.I(net15),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4546_ (.I(net16),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4547_ (.A1(_0433_),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4549_ (.A1(_0357_),
    .A2(_0431_),
    .B(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4550_ (.A1(net15),
    .A2(_3120_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4551_ (.I(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4552_ (.I(_0439_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4553_ (.I(\k.B[2][4] ),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4555_ (.A1(_0442_),
    .A2(_3312_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4556_ (.I(\k.B[2][3] ),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4557_ (.I(_0444_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4558_ (.A1(_3324_),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4559_ (.A1(_0443_),
    .A2(_0446_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4560_ (.A1(_0103_),
    .A2(_0445_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4561_ (.I(_0441_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4562_ (.I(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4563_ (.A1(_0450_),
    .A2(_3324_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4564_ (.A1(_0448_),
    .A2(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4565_ (.A1(_0452_),
    .A2(_0447_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4566_ (.I(\k.B[2][1] ),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4567_ (.A1(_0454_),
    .A2(_0070_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4568_ (.I(\k.B[2][0] ),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4569_ (.I(_0456_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4570_ (.I(_0457_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4571_ (.A1(_0458_),
    .A2(_0064_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4572_ (.I(\k.B[2][2] ),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4573_ (.I(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4574_ (.I(_0461_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4575_ (.A1(_3312_),
    .A2(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4576_ (.I(\k.B[2][1] ),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4577_ (.I(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4578_ (.I(_0465_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4579_ (.I(\k.B[2][0] ),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_0467_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4582_ (.A1(_0466_),
    .A2(_0064_),
    .B1(_0067_),
    .B2(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4583_ (.A1(_0455_),
    .A2(_0459_),
    .B1(_0463_),
    .B2(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_3330_),
    .A2(_0456_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4585_ (.A1(_0461_),
    .A2(_3315_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4586_ (.A1(_0472_),
    .A2(_0455_),
    .A3(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4587_ (.A1(_0471_),
    .A2(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(_0471_),
    .A2(_0474_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4589_ (.A1(_0453_),
    .A2(_0475_),
    .B(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4590_ (.I(\k.B[2][3] ),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4591_ (.A1(_3315_),
    .A2(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4592_ (.I(\k.B[2][5] ),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4593_ (.A1(_0480_),
    .A2(\k.A[3][0] ),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4594_ (.A1(_0479_),
    .A2(_0481_),
    .A3(_0443_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4595_ (.A1(_3329_),
    .A2(_0464_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4596_ (.A1(_0457_),
    .A2(_0067_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4597_ (.I(_0454_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4598_ (.A1(_0066_),
    .A2(_0457_),
    .B1(_0485_),
    .B2(_0067_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4599_ (.A1(_0483_),
    .A2(_0484_),
    .B1(_0473_),
    .B2(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4600_ (.A1(_0084_),
    .A2(_0467_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4601_ (.A1(_0460_),
    .A2(_3333_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4602_ (.A1(_0488_),
    .A2(_0483_),
    .A3(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4603_ (.A1(_0487_),
    .A2(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4604_ (.A1(_0482_),
    .A2(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4605_ (.A1(_0477_),
    .A2(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4606_ (.A1(_0447_),
    .A2(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4607_ (.A1(_0453_),
    .A2(_0475_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4608_ (.I(_0446_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4609_ (.I(_0485_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4610_ (.A1(_0497_),
    .A2(_0181_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4611_ (.I(_0469_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(_0499_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4613_ (.A1(_0500_),
    .A2(_0146_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4614_ (.I(_0461_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4615_ (.A1(_3325_),
    .A2(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4616_ (.I(_0466_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4617_ (.I(_0458_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4618_ (.A1(_0504_),
    .A2(_0195_),
    .B1(_0198_),
    .B2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4619_ (.A1(_0498_),
    .A2(_0501_),
    .B1(_0503_),
    .B2(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4620_ (.A1(_0484_),
    .A2(_0498_),
    .A3(_0463_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4621_ (.A1(_0507_),
    .A2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4622_ (.A1(_0507_),
    .A2(_0508_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4623_ (.A1(_0496_),
    .A2(_0509_),
    .B(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4624_ (.A1(_0495_),
    .A2(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4625_ (.A1(_0496_),
    .A2(_0509_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4626_ (.I(_0504_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4627_ (.A1(_0514_),
    .A2(_0146_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4628_ (.A1(_0459_),
    .A2(_0515_),
    .A3(_0503_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4629_ (.I(_0500_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4630_ (.A1(_0517_),
    .A2(_0127_),
    .A3(_0514_),
    .A4(_0256_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4631_ (.A1(_0516_),
    .A2(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4632_ (.A1(_0496_),
    .A2(_0509_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4633_ (.A1(_0513_),
    .A2(_0519_),
    .A3(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4634_ (.A1(_0512_),
    .A2(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4635_ (.A1(_0494_),
    .A2(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4636_ (.A1(_0477_),
    .A2(_0492_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4637_ (.A1(_0447_),
    .A2(_0493_),
    .B(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4638_ (.A1(_0441_),
    .A2(_3309_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4639_ (.A1(_0479_),
    .A2(_0443_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4640_ (.A1(_0526_),
    .A2(_0448_),
    .B1(_0527_),
    .B2(_0481_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4641_ (.I(\k.B[2][6] ),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4642_ (.I(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4643_ (.A1(_0530_),
    .A2(_0106_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4644_ (.A1(_0528_),
    .A2(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4645_ (.I(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4646_ (.A1(_0487_),
    .A2(_0490_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4647_ (.A1(_0482_),
    .A2(_0491_),
    .B(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4648_ (.A1(_0478_),
    .A2(_0070_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4649_ (.A1(_0480_),
    .A2(\k.A[3][1] ),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4650_ (.A1(_0536_),
    .A2(_0526_),
    .A3(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4651_ (.A1(_0072_),
    .A2(_0464_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4652_ (.A1(_0073_),
    .A2(_0456_),
    .B1(_0454_),
    .B2(_0086_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4653_ (.A1(_0539_),
    .A2(_0472_),
    .B1(_0489_),
    .B2(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4654_ (.A1(\k.A[3][4] ),
    .A2(_0460_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4655_ (.A1(_0090_),
    .A2(_0456_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4656_ (.A1(_0539_),
    .A2(_0542_),
    .A3(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4657_ (.A1(_0541_),
    .A2(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4658_ (.A1(_0538_),
    .A2(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4659_ (.A1(_0535_),
    .A2(_0546_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4660_ (.A1(_0533_),
    .A2(_0547_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4661_ (.A1(_0525_),
    .A2(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4662_ (.A1(_0495_),
    .A2(_0511_),
    .A3(_0494_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4663_ (.A1(_0549_),
    .A2(_0550_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4664_ (.A1(_0549_),
    .A2(_0550_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4665_ (.A1(_0523_),
    .A2(_0551_),
    .B(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4666_ (.A1(_0525_),
    .A2(_0548_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(_0530_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4668_ (.I(_0555_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4669_ (.I(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4670_ (.A1(_0557_),
    .A2(_0127_),
    .A3(_0528_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4671_ (.A1(_0535_),
    .A2(_0546_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4672_ (.A1(_0533_),
    .A2(_0547_),
    .B(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4673_ (.A1(_0536_),
    .A2(_0526_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4674_ (.A1(_0536_),
    .A2(_0526_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4675_ (.A1(_0537_),
    .A2(_0561_),
    .B(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4676_ (.A1(\k.B[2][6] ),
    .A2(_0103_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4677_ (.A1(\k.B[2][7] ),
    .A2(_3324_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4678_ (.A1(_0563_),
    .A2(_0564_),
    .A3(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4679_ (.A1(_0541_),
    .A2(_0544_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4680_ (.A1(_0538_),
    .A2(_0545_),
    .B(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4681_ (.A1(\k.B[2][4] ),
    .A2(_3332_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4682_ (.A1(\k.B[2][5] ),
    .A2(\k.A[3][2] ),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4683_ (.A1(_3330_),
    .A2(_0478_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4684_ (.A1(_0569_),
    .A2(_0570_),
    .A3(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4685_ (.A1(\k.A[3][6] ),
    .A2(\k.B[2][1] ),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4686_ (.A1(_0090_),
    .A2(_0467_),
    .B1(_0464_),
    .B2(_0084_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4687_ (.A1(_0488_),
    .A2(_0573_),
    .B1(_0574_),
    .B2(_0542_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4688_ (.A1(\k.A[3][5] ),
    .A2(\k.B[2][2] ),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4689_ (.A1(\k.A[3][7] ),
    .A2(_0467_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4690_ (.A1(_0573_),
    .A2(_0576_),
    .A3(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4691_ (.A1(_0575_),
    .A2(_0578_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4692_ (.A1(_0572_),
    .A2(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4693_ (.A1(_0568_),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4694_ (.A1(_0566_),
    .A2(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4695_ (.A1(_0560_),
    .A2(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4696_ (.A1(_0558_),
    .A2(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4697_ (.A1(_0554_),
    .A2(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4698_ (.A1(_0554_),
    .A2(_0584_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4699_ (.A1(_0553_),
    .A2(_0585_),
    .B(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4700_ (.A1(_0563_),
    .A2(_0564_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4701_ (.A1(_0563_),
    .A2(_0564_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4702_ (.A1(_0588_),
    .A2(_0565_),
    .B(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4703_ (.A1(_0568_),
    .A2(_0580_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4704_ (.A1(_0566_),
    .A2(_0581_),
    .B(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4705_ (.I(\k.B[2][7] ),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4706_ (.A1(_0593_),
    .A2(_0195_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4707_ (.A1(_0441_),
    .A2(_0086_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4708_ (.A1(_0569_),
    .A2(_0571_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4709_ (.A1(_0536_),
    .A2(_0595_),
    .B1(_0596_),
    .B2(_0570_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4710_ (.A1(_0529_),
    .A2(_0181_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4711_ (.A1(_0597_),
    .A2(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4712_ (.A1(_0594_),
    .A2(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4713_ (.A1(_0575_),
    .A2(_0578_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4714_ (.A1(_0572_),
    .A2(_0579_),
    .B(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4715_ (.A1(_0480_),
    .A2(_3333_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4716_ (.A1(_0153_),
    .A2(_0444_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4717_ (.A1(_0595_),
    .A2(_0603_),
    .A3(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4718_ (.A1(_0157_),
    .A2(_0468_),
    .B1(_0465_),
    .B2(_0160_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4719_ (.A1(_0157_),
    .A2(_0091_),
    .A3(_0468_),
    .A4(_0465_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4720_ (.A1(_0576_),
    .A2(_0606_),
    .B(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4721_ (.A1(_0157_),
    .A2(_0454_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4722_ (.A1(_0091_),
    .A2(_0460_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4723_ (.A1(_0609_),
    .A2(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4724_ (.A1(_0608_),
    .A2(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4725_ (.A1(_0605_),
    .A2(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4726_ (.A1(_0602_),
    .A2(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4727_ (.A1(_0600_),
    .A2(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4728_ (.A1(_0592_),
    .A2(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4729_ (.A1(_0590_),
    .A2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4730_ (.A1(_0533_),
    .A2(_0547_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4731_ (.A1(_0559_),
    .A2(_0618_),
    .B(_0582_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4732_ (.A1(_0558_),
    .A2(_0583_),
    .B(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4733_ (.I(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4734_ (.A1(_0617_),
    .A2(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4735_ (.A1(_0587_),
    .A2(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4736_ (.I(\k.B[0][4] ),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4737_ (.I(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(_0625_),
    .A2(_3129_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4739_ (.I(\k.B[0][3] ),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4740_ (.I(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4741_ (.A1(_0628_),
    .A2(_3137_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4742_ (.A1(_0626_),
    .A2(_0629_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4743_ (.A1(_0628_),
    .A2(_3130_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4744_ (.I(\k.B[0][4] ),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4745_ (.I(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4746_ (.A1(_0633_),
    .A2(_3189_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4747_ (.A1(_0631_),
    .A2(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4748_ (.A1(_0635_),
    .A2(_0630_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4749_ (.I(\k.B[0][1] ),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4750_ (.A1(_3144_),
    .A2(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4751_ (.I(\k.B[0][0] ),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4752_ (.I(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4753_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4754_ (.A1(_0641_),
    .A2(_3222_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4755_ (.I(\k.B[0][2] ),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4756_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4757_ (.A1(_3129_),
    .A2(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4758_ (.I(\k.B[0][1] ),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4759_ (.I(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4760_ (.I(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4761_ (.A1(_3145_),
    .A2(_0641_),
    .B1(_0648_),
    .B2(_3264_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4762_ (.A1(_0638_),
    .A2(_0642_),
    .B1(_0645_),
    .B2(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4763_ (.A1(_3142_),
    .A2(_0639_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4764_ (.I(_0643_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4765_ (.A1(_0652_),
    .A2(_3147_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4766_ (.A1(_0651_),
    .A2(_0638_),
    .A3(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4767_ (.A1(_0650_),
    .A2(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4768_ (.A1(_0650_),
    .A2(_0654_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4769_ (.A1(_0636_),
    .A2(_0655_),
    .B(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4770_ (.A1(_0627_),
    .A2(_3147_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4771_ (.I(\k.B[0][5] ),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4772_ (.A1(_0659_),
    .A2(\k.A[2][0] ),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4773_ (.A1(_0658_),
    .A2(_0660_),
    .A3(_0626_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4774_ (.A1(_3166_),
    .A2(_0646_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4775_ (.I(_0639_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4776_ (.A1(_3150_),
    .A2(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4777_ (.I(_0637_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4778_ (.A1(_3171_),
    .A2(_0640_),
    .B1(_0665_),
    .B2(_3150_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4779_ (.A1(_0662_),
    .A2(_0664_),
    .B1(_0653_),
    .B2(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4780_ (.I(\k.B[0][0] ),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4781_ (.A1(_3169_),
    .A2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4782_ (.A1(_3144_),
    .A2(_0652_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4783_ (.A1(_0669_),
    .A2(_0662_),
    .A3(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4784_ (.A1(_0667_),
    .A2(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4785_ (.A1(_0661_),
    .A2(_0672_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4786_ (.A1(_0657_),
    .A2(_0673_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4787_ (.A1(_0630_),
    .A2(_0675_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4788_ (.A1(_0636_),
    .A2(_0655_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4789_ (.I(_0629_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(_0648_),
    .A2(_3264_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4791_ (.I(_0640_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4792_ (.I(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4793_ (.A1(_0681_),
    .A2(_3276_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4794_ (.I(_0652_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4795_ (.A1(_3138_),
    .A2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4796_ (.I(_0665_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4797_ (.I(_0663_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4798_ (.A1(_0686_),
    .A2(_3276_),
    .B1(_3279_),
    .B2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4799_ (.A1(_0679_),
    .A2(_0682_),
    .B1(_0684_),
    .B2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4800_ (.A1(_0664_),
    .A2(_0679_),
    .A3(_0645_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4801_ (.A1(_0689_),
    .A2(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4802_ (.A1(_0689_),
    .A2(_0690_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4803_ (.A1(_0678_),
    .A2(_0691_),
    .B(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4804_ (.A1(_0677_),
    .A2(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4805_ (.A1(_0678_),
    .A2(_0691_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4806_ (.A1(_0686_),
    .A2(_3225_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4807_ (.A1(_0642_),
    .A2(_0697_),
    .A3(_0684_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4808_ (.I(_0681_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4809_ (.I(_0686_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4810_ (.A1(_0699_),
    .A2(_3207_),
    .A3(_0700_),
    .A4(_0252_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4811_ (.A1(_0698_),
    .A2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4812_ (.A1(_0678_),
    .A2(_0691_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4813_ (.A1(_0695_),
    .A2(_0702_),
    .A3(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4814_ (.A1(_0694_),
    .A2(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4815_ (.A1(_0676_),
    .A2(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4816_ (.A1(_0657_),
    .A2(_0673_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4817_ (.A1(_0630_),
    .A2(_0675_),
    .B(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4818_ (.A1(_0624_),
    .A2(_3126_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4819_ (.A1(_0658_),
    .A2(_0626_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4820_ (.A1(_0710_),
    .A2(_0631_),
    .B1(_0711_),
    .B2(_0660_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4821_ (.I(\k.B[0][6] ),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4822_ (.I(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4823_ (.A1(_0714_),
    .A2(_3138_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4824_ (.A1(_0712_),
    .A2(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4825_ (.I(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4826_ (.A1(_0667_),
    .A2(_0671_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4827_ (.A1(_0661_),
    .A2(_0672_),
    .B(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4828_ (.I(\k.B[0][3] ),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4829_ (.A1(_0721_),
    .A2(_3162_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4830_ (.A1(_0659_),
    .A2(\k.A[2][1] ),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4831_ (.A1(_0722_),
    .A2(_0710_),
    .A3(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4832_ (.A1(_3154_),
    .A2(_0646_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4833_ (.I(_0668_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4834_ (.I(_0646_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4835_ (.A1(_3155_),
    .A2(_0726_),
    .B1(_0727_),
    .B2(_3167_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4836_ (.A1(_0725_),
    .A2(_0651_),
    .B1(_0670_),
    .B2(_0728_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4837_ (.A1(_3166_),
    .A2(_0643_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4838_ (.A1(_3238_),
    .A2(_0639_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4839_ (.A1(_0725_),
    .A2(_0731_),
    .A3(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4840_ (.A1(_0730_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4841_ (.A1(_0724_),
    .A2(_0734_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4842_ (.A1(_0720_),
    .A2(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4843_ (.A1(_0717_),
    .A2(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4844_ (.A1(_0709_),
    .A2(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4845_ (.A1(_0677_),
    .A2(_0693_),
    .A3(_0676_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4846_ (.A1(_0738_),
    .A2(_0739_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4847_ (.A1(_0738_),
    .A2(_0739_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4848_ (.A1(_0706_),
    .A2(_0741_),
    .B(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4849_ (.A1(_0709_),
    .A2(_0737_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4850_ (.I(_0714_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4851_ (.I(_0745_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4852_ (.A1(_0746_),
    .A2(_3208_),
    .A3(_0712_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4853_ (.A1(_0720_),
    .A2(_0735_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4854_ (.A1(_0717_),
    .A2(_0736_),
    .B(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4855_ (.A1(_0722_),
    .A2(_0710_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4856_ (.A1(_0722_),
    .A2(_0710_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4857_ (.A1(_0723_),
    .A2(_0750_),
    .B(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4858_ (.A1(_0713_),
    .A2(_3187_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4859_ (.A1(\k.B[0][7] ),
    .A2(_3137_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4860_ (.A1(_0753_),
    .A2(_0754_),
    .A3(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4861_ (.A1(_0730_),
    .A2(_0733_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4862_ (.A1(_0724_),
    .A2(_0734_),
    .B(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4863_ (.A1(_0624_),
    .A2(_3162_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4864_ (.A1(\k.B[0][5] ),
    .A2(\k.A[2][2] ),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4865_ (.A1(_0721_),
    .A2(_3167_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4866_ (.A1(_0759_),
    .A2(_0760_),
    .A3(_0761_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4867_ (.A1(\k.A[2][6] ),
    .A2(\k.B[0][1] ),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4868_ (.A1(_3238_),
    .A2(_0668_),
    .B1(_0637_),
    .B2(_3169_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4869_ (.A1(_0669_),
    .A2(_0764_),
    .B1(_0765_),
    .B2(_0731_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4870_ (.A1(\k.A[2][5] ),
    .A2(\k.B[0][2] ),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4871_ (.A1(\k.A[2][7] ),
    .A2(_0668_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4872_ (.A1(_0764_),
    .A2(_0767_),
    .A3(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4873_ (.A1(_0766_),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4874_ (.A1(_0763_),
    .A2(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4875_ (.A1(_0758_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4876_ (.A1(_0756_),
    .A2(_0772_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4877_ (.A1(_0749_),
    .A2(_0774_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4878_ (.A1(_0747_),
    .A2(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4879_ (.A1(_0744_),
    .A2(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4880_ (.A1(_0744_),
    .A2(_0776_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4881_ (.A1(_0743_),
    .A2(_0777_),
    .B(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4882_ (.A1(_0753_),
    .A2(_0754_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4883_ (.A1(_0753_),
    .A2(_0754_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4884_ (.A1(_0780_),
    .A2(_0755_),
    .B(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4885_ (.A1(_0758_),
    .A2(_0771_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4886_ (.A1(_0756_),
    .A2(_0772_),
    .B(_0783_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4887_ (.I(\k.B[0][7] ),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4888_ (.A1(_0786_),
    .A2(_3225_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4889_ (.A1(_0624_),
    .A2(_3167_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4890_ (.A1(_0759_),
    .A2(_0761_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4891_ (.A1(_0722_),
    .A2(_0788_),
    .B1(_0789_),
    .B2(_0760_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4892_ (.A1(_0713_),
    .A2(_3279_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4893_ (.A1(_0790_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4894_ (.A1(_0787_),
    .A2(_0792_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4895_ (.A1(_0766_),
    .A2(_0769_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4896_ (.A1(_0763_),
    .A2(_0770_),
    .B(_0794_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4897_ (.A1(_0659_),
    .A2(_3150_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4898_ (.A1(_0627_),
    .A2(_3232_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4899_ (.A1(_0788_),
    .A2(_0797_),
    .A3(_0798_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4900_ (.A1(_3236_),
    .A2(_0726_),
    .B1(_0647_),
    .B2(_3175_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4901_ (.A1(_3236_),
    .A2(_3175_),
    .A3(_0726_),
    .A4(_0727_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4902_ (.A1(_0767_),
    .A2(_0800_),
    .B(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4903_ (.A1(\k.A[2][7] ),
    .A2(_0637_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_3238_),
    .A2(_0643_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4905_ (.A1(_0803_),
    .A2(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4906_ (.A1(_0802_),
    .A2(_0805_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4907_ (.A1(_0799_),
    .A2(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4908_ (.A1(_0796_),
    .A2(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4909_ (.A1(_0793_),
    .A2(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4910_ (.A1(_0785_),
    .A2(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4911_ (.A1(_0782_),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4912_ (.A1(_0717_),
    .A2(_0736_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4913_ (.A1(_0748_),
    .A2(_0813_),
    .B(_0774_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4914_ (.A1(_0747_),
    .A2(_0775_),
    .B(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4915_ (.I(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4916_ (.A1(_0812_),
    .A2(_0816_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4917_ (.A1(_0779_),
    .A2(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4918_ (.A1(_0623_),
    .A2(_0819_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4919_ (.A1(_0553_),
    .A2(_0585_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4920_ (.A1(_0743_),
    .A2(_0777_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4921_ (.A1(_0821_),
    .A2(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4922_ (.A1(_0523_),
    .A2(_0551_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4923_ (.A1(_0706_),
    .A2(_0741_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4924_ (.A1(_0824_),
    .A2(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4925_ (.A1(_0495_),
    .A2(_0511_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4926_ (.A1(_0512_),
    .A2(_0521_),
    .B(_0827_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4927_ (.A1(_0494_),
    .A2(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4928_ (.A1(_0677_),
    .A2(_0693_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4929_ (.A1(_0694_),
    .A2(_0704_),
    .B(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4930_ (.A1(_0676_),
    .A2(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4931_ (.A1(_0830_),
    .A2(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4932_ (.A1(_0512_),
    .A2(_0521_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4933_ (.A1(_0694_),
    .A2(_0704_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4934_ (.A1(_0835_),
    .A2(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4935_ (.A1(_0496_),
    .A2(_0509_),
    .A3(_0519_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4936_ (.A1(_0678_),
    .A2(_0691_),
    .A3(_0702_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4937_ (.A1(_0838_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4938_ (.A1(_0516_),
    .A2(_0518_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4939_ (.I(_0701_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4940_ (.A1(_0698_),
    .A2(_0843_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4941_ (.I(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4942_ (.A1(_0842_),
    .A2(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4943_ (.I(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4944_ (.I(_0514_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4945_ (.A1(_0127_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4946_ (.I(_0518_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4947_ (.A1(_0501_),
    .A2(_0849_),
    .B(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4948_ (.I(_0700_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4949_ (.A1(_3208_),
    .A2(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4950_ (.A1(_0682_),
    .A2(_0854_),
    .B(_0843_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4951_ (.A1(_0852_),
    .A2(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4952_ (.I(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4953_ (.A1(_0517_),
    .A2(_0699_),
    .A3(_3209_),
    .A4(_0128_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4954_ (.A1(_0852_),
    .A2(_0855_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4955_ (.A1(_0858_),
    .A2(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4956_ (.A1(_0842_),
    .A2(_0844_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4957_ (.I(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4958_ (.A1(_0857_),
    .A2(_0860_),
    .B(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4959_ (.A1(_0838_),
    .A2(_0840_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4960_ (.I(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4961_ (.A1(_0847_),
    .A2(_0864_),
    .B(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4962_ (.A1(_0835_),
    .A2(_0836_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4963_ (.A1(_0841_),
    .A2(_0867_),
    .B(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4964_ (.A1(_0830_),
    .A2(_0833_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4965_ (.A1(_0837_),
    .A2(_0869_),
    .B(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4966_ (.A1(_0834_),
    .A2(_0871_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4967_ (.A1(_0824_),
    .A2(_0825_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4968_ (.A1(_0826_),
    .A2(_0873_),
    .B(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4969_ (.A1(_0821_),
    .A2(_0822_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4970_ (.A1(_0823_),
    .A2(_0875_),
    .B(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4971_ (.A1(_0623_),
    .A2(_0819_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4972_ (.A1(_0820_),
    .A2(_0877_),
    .B(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4973_ (.A1(_0812_),
    .A2(_0816_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4974_ (.A1(_0779_),
    .A2(_0818_),
    .B(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4975_ (.I(_0746_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4976_ (.I(_0882_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4977_ (.A1(_0884_),
    .A2(_0403_),
    .A3(_0790_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4978_ (.I(_0786_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4979_ (.I(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4980_ (.I(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4981_ (.I(_0888_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4982_ (.A1(_0889_),
    .A2(_0252_),
    .A3(_0792_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4983_ (.A1(_0885_),
    .A2(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4984_ (.A1(_0796_),
    .A2(_0808_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4985_ (.A1(_0793_),
    .A2(_0809_),
    .B(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4986_ (.A1(_0786_),
    .A2(_0286_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4987_ (.A1(_0632_),
    .A2(_3232_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4988_ (.A1(_0788_),
    .A2(_0798_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4989_ (.A1(_0761_),
    .A2(_0896_),
    .B1(_0897_),
    .B2(_0797_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4990_ (.A1(_0714_),
    .A2(_3230_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4991_ (.A1(_0898_),
    .A2(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4992_ (.A1(_0895_),
    .A2(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4993_ (.A1(_0802_),
    .A2(_0805_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4994_ (.A1(_0799_),
    .A2(_0807_),
    .B(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4995_ (.I(_0659_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4996_ (.A1(_0904_),
    .A2(_3171_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4997_ (.A1(_0628_),
    .A2(_3243_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4998_ (.A1(_0896_),
    .A2(_0906_),
    .A3(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4999_ (.I(_0683_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5000_ (.A1(_3237_),
    .A2(_0909_),
    .A3(_0764_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5001_ (.A1(_0908_),
    .A2(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5002_ (.A1(_0903_),
    .A2(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5003_ (.A1(_0901_),
    .A2(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5004_ (.A1(_0893_),
    .A2(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5005_ (.A1(_0891_),
    .A2(_0914_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5006_ (.A1(_0891_),
    .A2(_0914_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5007_ (.A1(_0785_),
    .A2(_0810_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5008_ (.A1(_0782_),
    .A2(_0811_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5009_ (.A1(_0915_),
    .A2(_0917_),
    .B(_0918_),
    .C(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5010_ (.A1(_0918_),
    .A2(_0919_),
    .B(_0915_),
    .C(_0917_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5011_ (.I(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5012_ (.A1(_0920_),
    .A2(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5013_ (.A1(_0881_),
    .A2(_0923_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5014_ (.A1(_0617_),
    .A2(_0621_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5015_ (.A1(_0587_),
    .A2(_0622_),
    .B(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5016_ (.I(_0557_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5017_ (.A1(_0928_),
    .A2(_0323_),
    .A3(_0597_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5018_ (.I(_0593_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5019_ (.I(_0930_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5020_ (.I(_0931_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5021_ (.A1(_0932_),
    .A2(_0256_),
    .A3(_0599_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5022_ (.A1(_0929_),
    .A2(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5023_ (.A1(_0602_),
    .A2(_0613_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5024_ (.A1(_0600_),
    .A2(_0614_),
    .B(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5025_ (.A1(_0593_),
    .A2(_0143_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5026_ (.A1(_0449_),
    .A2(_0153_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5027_ (.A1(_0595_),
    .A2(_0604_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5028_ (.A1(_0571_),
    .A2(_0939_),
    .B1(_0940_),
    .B2(_0603_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5029_ (.A1(_0530_),
    .A2(_0334_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5030_ (.A1(_0937_),
    .A2(_0941_),
    .A3(_0942_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5031_ (.A1(_0608_),
    .A2(_0611_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5032_ (.A1(_0605_),
    .A2(_0612_),
    .B(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5033_ (.I(_0502_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5034_ (.A1(_0159_),
    .A2(_0946_),
    .A3(_0573_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5035_ (.I(_0480_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5036_ (.A1(_0948_),
    .A2(_0139_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5037_ (.A1(_0160_),
    .A2(_0444_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5038_ (.A1(_0939_),
    .A2(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5039_ (.A1(_0950_),
    .A2(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5040_ (.A1(_0947_),
    .A2(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5041_ (.A1(_0943_),
    .A2(_0945_),
    .A3(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5042_ (.A1(_0936_),
    .A2(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5043_ (.A1(_0934_),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5044_ (.A1(_0934_),
    .A2(_0956_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5045_ (.A1(_0592_),
    .A2(_0615_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5046_ (.A1(_0590_),
    .A2(_0616_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5047_ (.A1(_0957_),
    .A2(_0958_),
    .B(_0959_),
    .C(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5048_ (.A1(_0959_),
    .A2(_0961_),
    .B(_0957_),
    .C(_0958_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5049_ (.I(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5050_ (.A1(_0962_),
    .A2(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5051_ (.A1(_0926_),
    .A2(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5052_ (.A1(_0924_),
    .A2(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5053_ (.A1(_0924_),
    .A2(_0966_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5054_ (.A1(_0879_),
    .A2(_0967_),
    .B(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5055_ (.A1(_0936_),
    .A2(_0955_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5056_ (.A1(_0970_),
    .A2(_0957_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5057_ (.I(_0556_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5058_ (.A1(_0973_),
    .A2(_0362_),
    .B(_0941_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5059_ (.A1(_0973_),
    .A2(_0362_),
    .A3(_0941_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5060_ (.A1(_0937_),
    .A2(_0974_),
    .B(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5061_ (.A1(_0945_),
    .A2(_0954_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5062_ (.A1(_0945_),
    .A2(_0954_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5063_ (.A1(_0943_),
    .A2(_0977_),
    .B(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5064_ (.A1(_0930_),
    .A2(_0334_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5065_ (.A1(_0442_),
    .A2(_0161_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5066_ (.A1(_0604_),
    .A2(_0981_),
    .B1(_0952_),
    .B2(_0950_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5067_ (.A1(_0529_),
    .A2(_0375_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5068_ (.A1(_0983_),
    .A2(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5069_ (.A1(_0980_),
    .A2(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5070_ (.A1(_0609_),
    .A2(_0610_),
    .B1(_0947_),
    .B2(_0953_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5071_ (.I(_0948_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5072_ (.A1(_0988_),
    .A2(_0154_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5073_ (.I(_0478_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5074_ (.A1(_0158_),
    .A2(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5075_ (.A1(_0981_),
    .A2(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5076_ (.A1(_0989_),
    .A2(_0992_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5077_ (.A1(_0987_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5078_ (.A1(_0986_),
    .A2(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5079_ (.A1(_0979_),
    .A2(_0996_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5080_ (.A1(_0976_),
    .A2(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5081_ (.A1(_0972_),
    .A2(_0998_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5082_ (.A1(_0587_),
    .A2(_0622_),
    .B(_0964_),
    .C(_0925_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5083_ (.A1(_0962_),
    .A2(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5084_ (.A1(_0999_),
    .A2(_1001_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5085_ (.A1(_0893_),
    .A2(_0913_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5086_ (.A1(_1003_),
    .A2(_0915_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5087_ (.A1(_0882_),
    .A2(_0398_),
    .A3(_0898_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5088_ (.A1(_0888_),
    .A2(_0403_),
    .A3(_0900_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5089_ (.A1(_1006_),
    .A2(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5090_ (.A1(_0903_),
    .A2(_0911_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5091_ (.A1(_0901_),
    .A2(_0912_),
    .B(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5092_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0908_),
    .B2(_0910_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5093_ (.I(_0904_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5094_ (.A1(_1012_),
    .A2(_3233_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5095_ (.A1(_0625_),
    .A2(_3239_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5096_ (.I(_0721_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5097_ (.A1(_1016_),
    .A2(_3242_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5098_ (.A1(_1014_),
    .A2(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5099_ (.A1(_1013_),
    .A2(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5100_ (.A1(_1011_),
    .A2(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5101_ (.A1(_0786_),
    .A2(_0397_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5102_ (.A1(_0896_),
    .A2(_0907_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5103_ (.A1(_0798_),
    .A2(_1014_),
    .B1(_1022_),
    .B2(_0906_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5104_ (.A1(_0714_),
    .A2(_0412_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5105_ (.A1(_1023_),
    .A2(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5106_ (.A1(_1021_),
    .A2(_1025_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5107_ (.A1(_1020_),
    .A2(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5108_ (.A1(_1010_),
    .A2(_1028_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5109_ (.A1(_1008_),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5110_ (.A1(_1005_),
    .A2(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5111_ (.A1(_0779_),
    .A2(_0818_),
    .B(_0922_),
    .C(_0880_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5112_ (.A1(_0920_),
    .A2(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5113_ (.A1(_1031_),
    .A2(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5114_ (.A1(_1002_),
    .A2(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5115_ (.A1(_0969_),
    .A2(_1035_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5116_ (.A1(_0433_),
    .A2(net16),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5117_ (.I(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5118_ (.A1(_0432_),
    .A2(_0437_),
    .B1(_0440_),
    .B2(_1036_),
    .C(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5119_ (.I(net15),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5120_ (.A1(_1041_),
    .A2(_3120_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5121_ (.I(_1042_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5122_ (.A1(_0449_),
    .A2(_2754_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5123_ (.I(_0445_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5124_ (.A1(_2790_),
    .A2(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5125_ (.A1(_2755_),
    .A2(_0990_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5126_ (.A1(_0449_),
    .A2(_2740_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5127_ (.A1(_1047_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5128_ (.A1(_0988_),
    .A2(_2758_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5129_ (.A1(_1044_),
    .A2(_1046_),
    .B1(_1050_),
    .B2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5130_ (.A1(_0556_),
    .A2(_3001_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5131_ (.A1(_1052_),
    .A2(_1053_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5132_ (.A1(_1051_),
    .A2(_1050_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5133_ (.A1(_2821_),
    .A2(_0485_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5134_ (.A1(_2771_),
    .A2(_0499_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5135_ (.A1(_2755_),
    .A2(_0502_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5136_ (.A1(_2822_),
    .A2(_0458_),
    .B1(_0497_),
    .B2(_2771_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5137_ (.A1(_1056_),
    .A2(_1057_),
    .B1(_1058_),
    .B2(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5138_ (.A1(_2769_),
    .A2(_0461_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5139_ (.I(_2867_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5140_ (.A1(_1063_),
    .A2(_0469_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5141_ (.A1(_1056_),
    .A2(_1062_),
    .A3(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5142_ (.A1(_1061_),
    .A2(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5143_ (.A1(_1061_),
    .A2(_1065_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5144_ (.A1(_1055_),
    .A2(_1066_),
    .B(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5145_ (.A1(_0948_),
    .A2(_2740_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5146_ (.A1(_2769_),
    .A2(_0444_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5147_ (.A1(_1044_),
    .A2(_1069_),
    .A3(_1071_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5148_ (.I(_2811_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5149_ (.A1(_1073_),
    .A2(_0469_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5150_ (.A1(_2867_),
    .A2(_0465_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5151_ (.I(_1063_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5152_ (.A1(_1076_),
    .A2(_0458_),
    .B1(_0497_),
    .B2(_1073_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5153_ (.A1(_1074_),
    .A2(_1075_),
    .B1(_1077_),
    .B2(_1062_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5154_ (.A1(_2863_),
    .A2(_0468_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5155_ (.A1(_2821_),
    .A2(_0462_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5156_ (.A1(_1075_),
    .A2(_1079_),
    .A3(_1080_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5157_ (.A1(_1078_),
    .A2(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5158_ (.A1(_1072_),
    .A2(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5159_ (.A1(_1068_),
    .A2(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5160_ (.A1(_1068_),
    .A2(_1084_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5161_ (.A1(_1054_),
    .A2(_1085_),
    .B(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5162_ (.A1(_0593_),
    .A2(_3000_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5163_ (.A1(_2770_),
    .A2(_0442_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5164_ (.A1(_1044_),
    .A2(_1071_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5165_ (.A1(_1047_),
    .A2(_1089_),
    .B1(_1090_),
    .B2(_1069_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5166_ (.A1(_0529_),
    .A2(_2741_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5167_ (.A1(_1091_),
    .A2(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5168_ (.A1(_1088_),
    .A2(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5169_ (.A1(_1078_),
    .A2(_1082_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5170_ (.A1(_1072_),
    .A2(_1083_),
    .B(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5171_ (.I(_2862_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5172_ (.A1(_1098_),
    .A2(_0485_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5173_ (.I(_1098_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5174_ (.I(_0466_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5175_ (.A1(_1100_),
    .A2(_0499_),
    .B1(_1101_),
    .B2(_1076_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5176_ (.A1(_1064_),
    .A2(_1099_),
    .B1(_1102_),
    .B2(_1080_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5177_ (.A1(_2892_),
    .A2(_0457_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5178_ (.A1(_1063_),
    .A2(_0462_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5179_ (.A1(_1099_),
    .A2(_1105_),
    .A3(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5180_ (.A1(_1104_),
    .A2(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5181_ (.A1(_0988_),
    .A2(_2795_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5182_ (.A1(_1073_),
    .A2(_0990_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5183_ (.A1(_1089_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5184_ (.A1(_1109_),
    .A2(_1111_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5185_ (.A1(_1108_),
    .A2(_1112_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5186_ (.A1(_1095_),
    .A2(_1097_),
    .A3(_1113_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5187_ (.I(_3001_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5188_ (.A1(_0928_),
    .A2(_1116_),
    .A3(_1052_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5189_ (.A1(_1087_),
    .A2(_1115_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5190_ (.A1(_1117_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5191_ (.A1(_1087_),
    .A2(_1115_),
    .B(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5192_ (.I(_0928_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5193_ (.I(_3005_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5194_ (.A1(_1121_),
    .A2(_1122_),
    .A3(_1091_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5195_ (.I(_0932_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5196_ (.I(_1116_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5197_ (.A1(_1124_),
    .A2(_1126_),
    .A3(_1094_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5198_ (.A1(_1123_),
    .A2(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5199_ (.A1(_1097_),
    .A2(_1113_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5200_ (.A1(_1097_),
    .A2(_1113_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5201_ (.A1(_1095_),
    .A2(_1129_),
    .B(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5202_ (.A1(_1104_),
    .A2(_1107_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5203_ (.A1(_1108_),
    .A2(_1112_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5204_ (.A1(_1132_),
    .A2(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5205_ (.I(_2770_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5206_ (.A1(_1135_),
    .A2(_0988_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5207_ (.A1(_1073_),
    .A2(_0450_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5208_ (.A1(_1063_),
    .A2(_0445_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5209_ (.A1(_1138_),
    .A2(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5210_ (.A1(_1137_),
    .A2(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5211_ (.A1(_2892_),
    .A2(_0497_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5212_ (.A1(_1098_),
    .A2(_0462_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5213_ (.A1(_1142_),
    .A2(_1143_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5214_ (.A1(_2926_),
    .A2(_0505_),
    .B1(_1101_),
    .B2(_1100_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5215_ (.A1(_1100_),
    .A2(_2926_),
    .A3(_0499_),
    .A4(_1101_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5216_ (.A1(_1145_),
    .A2(_1106_),
    .B(_1146_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5217_ (.A1(_1144_),
    .A2(_1148_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5218_ (.A1(_1141_),
    .A2(_1149_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5219_ (.A1(_1134_),
    .A2(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5220_ (.A1(_0930_),
    .A2(_3005_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5221_ (.A1(_1071_),
    .A2(_1138_),
    .B1(_1111_),
    .B2(_1109_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5222_ (.A1(_0530_),
    .A2(_2792_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5223_ (.A1(_1153_),
    .A2(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5224_ (.A1(_1152_),
    .A2(_1155_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5225_ (.I(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5226_ (.A1(_1151_),
    .A2(_1157_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5227_ (.A1(_1131_),
    .A2(_1159_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5228_ (.A1(_1128_),
    .A2(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5229_ (.A1(_2758_),
    .A2(_1045_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5230_ (.A1(_1049_),
    .A2(_1162_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5231_ (.I(_0450_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5232_ (.A1(_1164_),
    .A2(_3000_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5233_ (.A1(_1046_),
    .A2(_1165_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5234_ (.A1(_1166_),
    .A2(_1163_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5235_ (.A1(_2770_),
    .A2(_0466_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5236_ (.A1(_0505_),
    .A2(_2795_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5237_ (.A1(_2741_),
    .A2(_0502_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5238_ (.A1(_1135_),
    .A2(_0505_),
    .B1(_0504_),
    .B2(_2795_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5239_ (.A1(_1168_),
    .A2(_1170_),
    .B1(_1171_),
    .B2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5240_ (.A1(_1074_),
    .A2(_1168_),
    .A3(_1058_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5241_ (.A1(_1173_),
    .A2(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5242_ (.A1(_1173_),
    .A2(_1174_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5243_ (.A1(_1167_),
    .A2(_1175_),
    .B(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5244_ (.A1(_1055_),
    .A2(_1066_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5245_ (.A1(_1177_),
    .A2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5246_ (.A1(_1163_),
    .A2(_1179_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5247_ (.A1(_1167_),
    .A2(_1175_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5248_ (.A1(_1101_),
    .A2(_2778_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5249_ (.A1(_0500_),
    .A2(_3002_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5250_ (.A1(_3002_),
    .A2(_0504_),
    .B1(_2792_),
    .B2(_0500_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5251_ (.A1(_3000_),
    .A2(_0946_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5252_ (.A1(_1183_),
    .A2(_1184_),
    .B1(_1185_),
    .B2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5253_ (.A1(_1057_),
    .A2(_1183_),
    .A3(_1171_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5254_ (.A1(_1187_),
    .A2(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5255_ (.A1(_1187_),
    .A2(_1188_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5256_ (.A1(_1162_),
    .A2(_1189_),
    .B(_1190_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5257_ (.A1(_1182_),
    .A2(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5258_ (.A1(_3005_),
    .A2(_0514_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5259_ (.A1(_1170_),
    .A2(_1194_),
    .A3(_1186_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5260_ (.A1(_1116_),
    .A2(_0517_),
    .A3(_1122_),
    .A4(_0848_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5261_ (.A1(_1162_),
    .A2(_1189_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5262_ (.A1(_1195_),
    .A2(_1196_),
    .A3(_1197_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5263_ (.A1(_1181_),
    .A2(_1193_),
    .A3(_1198_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5264_ (.A1(_1068_),
    .A2(_1084_),
    .A3(_1054_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5265_ (.A1(_1177_),
    .A2(_1178_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5266_ (.A1(_1163_),
    .A2(_1179_),
    .B(_1201_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5267_ (.A1(_1200_),
    .A2(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5268_ (.A1(_1182_),
    .A2(_1192_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5269_ (.A1(_1205_),
    .A2(_1181_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5270_ (.A1(_1204_),
    .A2(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5271_ (.A1(_1204_),
    .A2(_1206_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5272_ (.A1(_1199_),
    .A2(_1207_),
    .B(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5273_ (.A1(_1200_),
    .A2(_1203_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5274_ (.A1(_1117_),
    .A2(_1118_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5275_ (.A1(_1210_),
    .A2(_1211_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5276_ (.A1(_1210_),
    .A2(_1211_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5277_ (.A1(_1209_),
    .A2(_1212_),
    .B(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5278_ (.A1(_1120_),
    .A2(_1161_),
    .A3(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5279_ (.A1(_0632_),
    .A2(_0927_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5280_ (.I(_0628_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5281_ (.A1(_1218_),
    .A2(_2499_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5282_ (.A1(_0627_),
    .A2(_0938_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5283_ (.A1(_0632_),
    .A2(_0960_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5284_ (.A1(_1220_),
    .A2(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5285_ (.A1(_1012_),
    .A2(_0806_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5286_ (.A1(_1217_),
    .A2(_1219_),
    .B1(_1222_),
    .B2(_1223_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5287_ (.A1(_0745_),
    .A2(_2102_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5288_ (.A1(_1225_),
    .A2(_1226_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5289_ (.A1(_1223_),
    .A2(_1222_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5290_ (.A1(_1290_),
    .A2(_0727_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5291_ (.A1(_2719_),
    .A2(_0680_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5292_ (.A1(_1433_),
    .A2(_0683_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5293_ (.A1(_3110_),
    .A2(_0641_),
    .B1(_0648_),
    .B2(_2719_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5294_ (.A1(_1229_),
    .A2(_1230_),
    .B1(_1231_),
    .B2(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5295_ (.A1(_1257_),
    .A2(_0652_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5296_ (.A1(_3099_),
    .A2(_0663_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5297_ (.A1(_1229_),
    .A2(_1234_),
    .A3(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5298_ (.A1(_1233_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5299_ (.A1(_1233_),
    .A2(_1237_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5300_ (.A1(_1228_),
    .A2(_1238_),
    .B(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5301_ (.A1(_0904_),
    .A2(_0762_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5302_ (.A1(_0721_),
    .A2(_1257_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5303_ (.A1(_1217_),
    .A2(_1241_),
    .A3(_1242_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5304_ (.I(_1290_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5305_ (.A1(_1244_),
    .A2(_0663_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5306_ (.A1(_3099_),
    .A2(_0727_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5307_ (.I(_3099_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5308_ (.A1(_1248_),
    .A2(_0641_),
    .B1(_0665_),
    .B2(_1244_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5309_ (.A1(_1245_),
    .A2(_1247_),
    .B1(_1249_),
    .B2(_1234_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5310_ (.A1(_2298_),
    .A2(_0726_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5311_ (.A1(_1244_),
    .A2(_0644_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5312_ (.A1(_1247_),
    .A2(_1251_),
    .A3(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5313_ (.A1(_1250_),
    .A2(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5314_ (.A1(_1243_),
    .A2(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5315_ (.A1(_1240_),
    .A2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5316_ (.A1(_1240_),
    .A2(_1255_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5317_ (.A1(_1227_),
    .A2(_1256_),
    .B(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5318_ (.A1(\k.B[0][7] ),
    .A2(_1652_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5319_ (.A1(_0625_),
    .A2(_1015_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5320_ (.A1(_1217_),
    .A2(_1242_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5321_ (.A1(_1220_),
    .A2(_1261_),
    .B1(_1262_),
    .B2(_1241_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5322_ (.A1(\k.B[0][6] ),
    .A2(_0762_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5323_ (.A1(_1263_),
    .A2(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5324_ (.A1(_1260_),
    .A2(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5325_ (.A1(_1250_),
    .A2(_1253_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5326_ (.A1(_1243_),
    .A2(_1254_),
    .B(_1267_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5327_ (.A1(_2726_),
    .A2(_0647_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5328_ (.I(_2726_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5329_ (.I(_0647_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5330_ (.A1(_1271_),
    .A2(_0680_),
    .B1(_1272_),
    .B2(_3100_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5331_ (.A1(_1236_),
    .A2(_1270_),
    .B1(_1273_),
    .B2(_1252_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5332_ (.A1(_2671_),
    .A2(_0640_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5333_ (.A1(_1248_),
    .A2(_0644_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5334_ (.A1(_1270_),
    .A2(_1275_),
    .A3(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5335_ (.A1(_1274_),
    .A2(_1277_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5336_ (.A1(_1012_),
    .A2(_2705_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5337_ (.A1(_1016_),
    .A2(_1244_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5338_ (.A1(_1261_),
    .A2(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5339_ (.A1(_1280_),
    .A2(_1282_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5340_ (.A1(_1278_),
    .A2(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5341_ (.A1(_1266_),
    .A2(_1269_),
    .A3(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5342_ (.I(_2102_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5343_ (.A1(_0884_),
    .A2(_1286_),
    .A3(_1225_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5344_ (.A1(_1259_),
    .A2(_1285_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5345_ (.A1(_1287_),
    .A2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5346_ (.A1(_1259_),
    .A2(_1285_),
    .B(_1289_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5347_ (.I(_0884_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5348_ (.A1(_1292_),
    .A2(_2710_),
    .A3(_1263_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5349_ (.I(_0889_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5350_ (.I(_1286_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5351_ (.A1(_1294_),
    .A2(_1295_),
    .A3(_1265_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5352_ (.A1(_1293_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5353_ (.A1(_1269_),
    .A2(_1284_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5354_ (.A1(_1269_),
    .A2(_1284_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5355_ (.A1(_1266_),
    .A2(_1298_),
    .B(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5356_ (.A1(_1274_),
    .A2(_1277_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5357_ (.A1(_1278_),
    .A2(_1283_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5358_ (.A1(_1302_),
    .A2(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5359_ (.A1(_1012_),
    .A2(_3089_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5360_ (.A1(_0633_),
    .A2(_3110_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5361_ (.A1(_1016_),
    .A2(_1248_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5362_ (.A1(_1306_),
    .A2(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5363_ (.A1(_1305_),
    .A2(_1308_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5364_ (.A1(_2729_),
    .A2(_0648_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5365_ (.A1(_1271_),
    .A2(_0644_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5366_ (.A1(_1310_),
    .A2(_1311_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5367_ (.I(_1271_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5368_ (.A1(_2729_),
    .A2(_0687_),
    .B1(_1272_),
    .B2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5369_ (.I(_2729_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5370_ (.A1(_1316_),
    .A2(_1314_),
    .A3(_0680_),
    .A4(_1272_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5371_ (.A1(_1315_),
    .A2(_1276_),
    .B(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5372_ (.A1(_1313_),
    .A2(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5373_ (.A1(_1309_),
    .A2(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5374_ (.A1(_1304_),
    .A2(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5375_ (.A1(_0886_),
    .A2(_2519_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5376_ (.A1(_1242_),
    .A2(_1306_),
    .B1(_1282_),
    .B2(_1280_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5377_ (.I(_0713_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5378_ (.A1(_1325_),
    .A2(_2705_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5379_ (.A1(_1324_),
    .A2(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5380_ (.A1(_1322_),
    .A2(_1327_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5381_ (.I(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5382_ (.A1(_1321_),
    .A2(_1329_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5383_ (.A1(_1300_),
    .A2(_1330_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5384_ (.A1(_1297_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5385_ (.A1(_1218_),
    .A2(_1652_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5386_ (.A1(_1221_),
    .A2(_1333_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5387_ (.I(_0633_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5388_ (.A1(_1336_),
    .A2(_1652_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5389_ (.A1(_1219_),
    .A2(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5390_ (.A1(_1338_),
    .A2(_1335_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5391_ (.A1(_1015_),
    .A2(_0665_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5392_ (.A1(_0687_),
    .A2(_1521_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5393_ (.A1(_1466_),
    .A2(_0683_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5394_ (.A1(_3089_),
    .A2(_0687_),
    .B1(_0686_),
    .B2(_1521_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5395_ (.A1(_1340_),
    .A2(_1341_),
    .B1(_1342_),
    .B2(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5396_ (.A1(_1245_),
    .A2(_1340_),
    .A3(_1231_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5397_ (.A1(_1344_),
    .A2(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5398_ (.A1(_1344_),
    .A2(_1346_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5399_ (.A1(_1339_),
    .A2(_1347_),
    .B(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5400_ (.A1(_1228_),
    .A2(_1238_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5401_ (.A1(_1349_),
    .A2(_1350_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5402_ (.A1(_1335_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5403_ (.A1(_1339_),
    .A2(_1347_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5404_ (.A1(_1272_),
    .A2(_1521_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5405_ (.A1(_0681_),
    .A2(_2509_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5406_ (.A1(_2499_),
    .A2(_0700_),
    .B1(_2706_),
    .B2(_0681_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5407_ (.A1(_1663_),
    .A2(_0909_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5408_ (.A1(_1354_),
    .A2(_1355_),
    .B1(_1357_),
    .B2(_1358_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5409_ (.A1(_1230_),
    .A2(_1354_),
    .A3(_1342_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5410_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5411_ (.A1(_1359_),
    .A2(_1360_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5412_ (.A1(_1333_),
    .A2(_1361_),
    .B(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5413_ (.A1(_1353_),
    .A2(_1363_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5414_ (.A1(_1333_),
    .A2(_1361_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5415_ (.A1(_2509_),
    .A2(_0700_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5416_ (.A1(_1341_),
    .A2(_1366_),
    .A3(_1358_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5417_ (.A1(_0699_),
    .A2(_1286_),
    .A3(_2519_),
    .A4(_0853_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5418_ (.A1(_1368_),
    .A2(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5419_ (.A1(_1333_),
    .A2(_1361_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5420_ (.A1(_1365_),
    .A2(_1370_),
    .A3(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5421_ (.I(_1372_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5422_ (.A1(_1352_),
    .A2(_1364_),
    .A3(_1373_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5423_ (.A1(_1240_),
    .A2(_1255_),
    .A3(_1227_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5424_ (.A1(_1349_),
    .A2(_1350_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5425_ (.A1(_1335_),
    .A2(_1351_),
    .B(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5426_ (.A1(_1375_),
    .A2(_1377_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5427_ (.A1(_1353_),
    .A2(_1363_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5428_ (.A1(_1380_),
    .A2(_1352_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5429_ (.A1(_1379_),
    .A2(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5430_ (.A1(_1379_),
    .A2(_1381_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5431_ (.A1(_1374_),
    .A2(_1382_),
    .B(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5432_ (.A1(_1375_),
    .A2(_1377_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5433_ (.A1(_1287_),
    .A2(_1288_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5434_ (.A1(_1385_),
    .A2(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5435_ (.A1(_1385_),
    .A2(_1386_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5436_ (.A1(_1384_),
    .A2(_1387_),
    .B(_1388_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5437_ (.A1(_1291_),
    .A2(_1332_),
    .A3(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5438_ (.A1(_1216_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5439_ (.A1(_1181_),
    .A2(_1193_),
    .A3(_1198_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5440_ (.A1(_1204_),
    .A2(_1206_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5441_ (.A1(_1204_),
    .A2(_1206_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5442_ (.A1(_1393_),
    .A2(_1394_),
    .B(_1395_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5443_ (.A1(_1396_),
    .A2(_1212_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5444_ (.A1(_1352_),
    .A2(_1364_),
    .A3(_1373_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5445_ (.A1(_1379_),
    .A2(_1381_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5446_ (.A1(_1379_),
    .A2(_1381_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5447_ (.A1(_1398_),
    .A2(_1399_),
    .B(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5448_ (.A1(_1402_),
    .A2(_1387_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5449_ (.A1(_1397_),
    .A2(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5450_ (.A1(_1393_),
    .A2(_1394_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5451_ (.A1(_1199_),
    .A2(_1207_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5452_ (.A1(_1374_),
    .A2(_1382_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5453_ (.A1(_1398_),
    .A2(_1399_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5454_ (.A1(_1405_),
    .A2(_1406_),
    .B1(_1407_),
    .B2(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5455_ (.A1(_1193_),
    .A2(_1198_),
    .B(_1205_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5456_ (.A1(_1181_),
    .A2(_1410_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5457_ (.A1(_1364_),
    .A2(_1373_),
    .B(_1380_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5458_ (.A1(_1352_),
    .A2(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5459_ (.A1(_1412_),
    .A2(_1414_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5460_ (.A1(_1193_),
    .A2(_1198_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5461_ (.A1(_1364_),
    .A2(_1372_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5462_ (.A1(_1416_),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5463_ (.A1(_1195_),
    .A2(_1196_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5464_ (.A1(_1419_),
    .A2(_1197_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5465_ (.A1(_1365_),
    .A2(_1371_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5466_ (.A1(_1368_),
    .A2(_1369_),
    .B(_1421_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5467_ (.A1(_1373_),
    .A2(_1420_),
    .A3(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5468_ (.A1(_1370_),
    .A2(_1421_),
    .A3(_1420_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5469_ (.A1(_1116_),
    .A2(_0848_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5470_ (.A1(_1184_),
    .A2(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5471_ (.A1(_1196_),
    .A2(_1427_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5472_ (.A1(_1286_),
    .A2(_0853_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5473_ (.A1(_1355_),
    .A2(_1429_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5474_ (.A1(_1369_),
    .A2(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5475_ (.A1(_1428_),
    .A2(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5476_ (.I(_0517_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5477_ (.I(_0699_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5478_ (.A1(_1126_),
    .A2(_1434_),
    .A3(_1435_),
    .A4(_1295_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5479_ (.A1(_1428_),
    .A2(_1431_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5480_ (.A1(_1432_),
    .A2(_1436_),
    .B(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5481_ (.A1(_1195_),
    .A2(_1196_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5482_ (.A1(_1368_),
    .A2(_1369_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5483_ (.A1(_1439_),
    .A2(_1440_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5484_ (.A1(_1439_),
    .A2(_1440_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5485_ (.A1(_1438_),
    .A2(_1441_),
    .B(_1442_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5486_ (.A1(_1425_),
    .A2(_1443_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5487_ (.A1(_1416_),
    .A2(_1417_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5488_ (.A1(_1424_),
    .A2(_1445_),
    .B(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5489_ (.A1(_1412_),
    .A2(_1414_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5490_ (.A1(_1418_),
    .A2(_1447_),
    .B(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5491_ (.A1(_1415_),
    .A2(_1449_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5492_ (.A1(_1405_),
    .A2(_1408_),
    .A3(_1406_),
    .A4(_1407_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5493_ (.A1(_1409_),
    .A2(_1450_),
    .B(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5494_ (.A1(_1397_),
    .A2(_1403_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5495_ (.A1(_1404_),
    .A2(_1452_),
    .B(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5496_ (.A1(_1216_),
    .A2(_1391_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5497_ (.A1(_1392_),
    .A2(_1454_),
    .B(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5498_ (.A1(_1120_),
    .A2(_1161_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5499_ (.A1(_1120_),
    .A2(_1161_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5500_ (.A1(_1215_),
    .A2(_1458_),
    .B(_1459_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5501_ (.A1(_1131_),
    .A2(_1159_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5502_ (.A1(_1128_),
    .A2(_1160_),
    .B(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5503_ (.I(_2792_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5504_ (.A1(_1121_),
    .A2(_1463_),
    .A3(_1153_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5505_ (.I(_1124_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5506_ (.A1(_1465_),
    .A2(_1122_),
    .A3(_1155_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5507_ (.A1(_1464_),
    .A2(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5508_ (.A1(_1134_),
    .A2(_1150_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5509_ (.A1(_1151_),
    .A2(_1157_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5510_ (.A1(_1469_),
    .A2(_1470_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5511_ (.A1(_1144_),
    .A2(_1148_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5512_ (.A1(_1141_),
    .A2(_1149_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5513_ (.A1(_1472_),
    .A2(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5514_ (.A1(_2956_),
    .A2(_0946_),
    .A3(_1099_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5515_ (.I(_0948_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5516_ (.A1(_2822_),
    .A2(_1476_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5517_ (.A1(_1076_),
    .A2(_0442_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5518_ (.A1(_1098_),
    .A2(_0990_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5519_ (.A1(_1479_),
    .A2(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5520_ (.A1(_1478_),
    .A2(_1481_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5521_ (.A1(_1475_),
    .A2(_1482_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5522_ (.A1(_1474_),
    .A2(_1483_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5523_ (.A1(_0930_),
    .A2(_1463_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5524_ (.A1(_1110_),
    .A2(_1479_),
    .B1(_1140_),
    .B2(_1137_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5525_ (.A1(_1135_),
    .A2(_0555_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5526_ (.A1(_1486_),
    .A2(_1487_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5527_ (.A1(_1485_),
    .A2(_1489_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5528_ (.I(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5529_ (.A1(_1484_),
    .A2(_1491_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5530_ (.A1(_1471_),
    .A2(_1492_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5531_ (.A1(_1468_),
    .A2(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5532_ (.A1(_1462_),
    .A2(_1494_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5533_ (.A1(_1460_),
    .A2(_1495_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5534_ (.A1(_1291_),
    .A2(_1332_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5535_ (.A1(_1291_),
    .A2(_1332_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5536_ (.A1(_1390_),
    .A2(_1497_),
    .B(_1498_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5537_ (.A1(_1300_),
    .A2(_1330_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5538_ (.A1(_1297_),
    .A2(_1331_),
    .B(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5539_ (.A1(_1292_),
    .A2(_3092_),
    .A3(_1324_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5540_ (.A1(_1294_),
    .A2(_2710_),
    .A3(_1327_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5541_ (.A1(_1503_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5542_ (.A1(_1304_),
    .A2(_1320_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5543_ (.A1(_1321_),
    .A2(_1329_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5544_ (.A1(_1506_),
    .A2(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5545_ (.A1(_1313_),
    .A2(_1318_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5546_ (.A1(_1309_),
    .A2(_1319_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5547_ (.A1(_1509_),
    .A2(_1511_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5548_ (.I(_1316_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5549_ (.A1(_1513_),
    .A2(_0909_),
    .A3(_1270_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5550_ (.I(_0904_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5551_ (.I(_3110_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5552_ (.A1(_1515_),
    .A2(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5553_ (.A1(_0625_),
    .A2(_1248_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5554_ (.A1(_1016_),
    .A2(_1271_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5555_ (.A1(_1518_),
    .A2(_1519_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5556_ (.A1(_1517_),
    .A2(_1520_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5557_ (.A1(_1514_),
    .A2(_1522_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5558_ (.A1(_1512_),
    .A2(_1523_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5559_ (.A1(_0886_),
    .A2(_2706_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5560_ (.A1(_1281_),
    .A2(_1518_),
    .B1(_1308_),
    .B2(_1305_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5561_ (.A1(_1325_),
    .A2(_3090_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5562_ (.A1(_1526_),
    .A2(_1527_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5563_ (.A1(_1525_),
    .A2(_1528_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5564_ (.I(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5565_ (.A1(_1524_),
    .A2(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5566_ (.A1(_1508_),
    .A2(_1531_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5567_ (.A1(_1505_),
    .A2(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5568_ (.A1(_1502_),
    .A2(_1534_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5569_ (.A1(_1500_),
    .A2(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5570_ (.A1(_1496_),
    .A2(_1536_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5571_ (.A1(_1496_),
    .A2(_1536_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5572_ (.A1(_1457_),
    .A2(_1537_),
    .B(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5573_ (.A1(_1502_),
    .A2(_1534_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5574_ (.A1(_1500_),
    .A2(_1535_),
    .B(_1540_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5575_ (.A1(_1508_),
    .A2(_1531_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5576_ (.A1(_1505_),
    .A2(_1533_),
    .B(_1542_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5577_ (.I(_0884_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5578_ (.I(_3090_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5579_ (.A1(_1545_),
    .A2(_1546_),
    .A3(_1526_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5580_ (.I(_0889_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5581_ (.A1(_1548_),
    .A2(_3092_),
    .A3(_1528_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5582_ (.A1(_1547_),
    .A2(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5583_ (.A1(_1512_),
    .A2(_1523_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5584_ (.A1(_1524_),
    .A2(_1530_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5585_ (.A1(_1551_),
    .A2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5586_ (.A1(_0887_),
    .A2(_3090_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5587_ (.A1(_0633_),
    .A2(_1314_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5588_ (.A1(_1307_),
    .A2(_1556_),
    .B1(_1520_),
    .B2(_1517_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5589_ (.A1(_1325_),
    .A2(_1516_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5590_ (.A1(_1557_),
    .A2(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5591_ (.A1(_1555_),
    .A2(_1559_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5592_ (.A1(_1310_),
    .A2(_1311_),
    .B1(_1514_),
    .B2(_1522_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5593_ (.I(_3100_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5594_ (.A1(_1515_),
    .A2(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5595_ (.A1(_1218_),
    .A2(_1316_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5596_ (.A1(_1556_),
    .A2(_1564_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5597_ (.A1(_1563_),
    .A2(_1566_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5598_ (.A1(_1561_),
    .A2(_1567_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5599_ (.A1(_1560_),
    .A2(_1568_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5600_ (.A1(_1553_),
    .A2(_1569_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5601_ (.A1(_1550_),
    .A2(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5602_ (.A1(_1544_),
    .A2(_1571_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5603_ (.A1(_1541_),
    .A2(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5604_ (.A1(_1462_),
    .A2(_1494_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5605_ (.A1(_1460_),
    .A2(_1495_),
    .B(_1574_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5606_ (.A1(_1471_),
    .A2(_1492_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5607_ (.A1(_1468_),
    .A2(_1493_),
    .B(_1577_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5608_ (.I(_1135_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5609_ (.I(_0928_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5610_ (.A1(_1579_),
    .A2(_1580_),
    .A3(_1486_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5611_ (.I(_1124_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5612_ (.A1(_1582_),
    .A2(_1463_),
    .A3(_1489_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5613_ (.A1(_1581_),
    .A2(_1583_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5614_ (.A1(_1474_),
    .A2(_1483_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5615_ (.A1(_1484_),
    .A2(_1491_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5616_ (.A1(_1585_),
    .A2(_1586_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5617_ (.A1(_1579_),
    .A2(_0931_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5618_ (.I(_1100_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5619_ (.A1(_1590_),
    .A2(_0450_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5620_ (.A1(_1139_),
    .A2(_1591_),
    .B1(_1481_),
    .B2(_1478_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5621_ (.I(_2822_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5622_ (.A1(_1593_),
    .A2(_0555_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5623_ (.A1(_1592_),
    .A2(_1594_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5624_ (.A1(_1589_),
    .A2(_1595_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5625_ (.A1(_1142_),
    .A2(_1143_),
    .B1(_1475_),
    .B2(_1482_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5626_ (.I(_1076_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5627_ (.A1(_1599_),
    .A2(_1476_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5628_ (.A1(_2956_),
    .A2(_1045_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5629_ (.A1(_1591_),
    .A2(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5630_ (.A1(_1600_),
    .A2(_1602_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5631_ (.A1(_1597_),
    .A2(_1603_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5632_ (.A1(_1596_),
    .A2(_1604_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5633_ (.A1(_1588_),
    .A2(_1605_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5634_ (.A1(_1584_),
    .A2(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5635_ (.A1(_1578_),
    .A2(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5636_ (.A1(_1575_),
    .A2(_1608_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5637_ (.A1(_1539_),
    .A2(_1573_),
    .A3(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5638_ (.A1(_1043_),
    .A2(_1611_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5639_ (.I(net1),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5640_ (.I(_1613_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5641_ (.A1(_3125_),
    .A2(_1040_),
    .B(_1612_),
    .C(_1614_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5642_ (.I(_1038_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5643_ (.I(_1615_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5644_ (.I(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5645_ (.A1(_1573_),
    .A2(_1610_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5646_ (.A1(_1573_),
    .A2(_1610_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5647_ (.A1(_1539_),
    .A2(_1618_),
    .B(_1620_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5648_ (.A1(_1544_),
    .A2(_1571_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5649_ (.A1(_1541_),
    .A2(_1572_),
    .B(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5650_ (.A1(_1553_),
    .A2(_1569_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5651_ (.A1(_1550_),
    .A2(_1570_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5652_ (.A1(_1624_),
    .A2(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5653_ (.I(_1516_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5654_ (.A1(_1292_),
    .A2(_1627_),
    .A3(_1557_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5655_ (.A1(_1294_),
    .A2(_1546_),
    .A3(_1559_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5656_ (.A1(_1628_),
    .A2(_1629_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(_1336_),
    .A2(_1513_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5658_ (.I(_1515_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5659_ (.I(_1314_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5660_ (.I(_1634_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5661_ (.A1(_1633_),
    .A2(_1635_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5662_ (.I(_1513_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5663_ (.A1(_1633_),
    .A2(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5664_ (.A1(_1556_),
    .A2(_1638_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5665_ (.A1(_1632_),
    .A2(_1636_),
    .B(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5666_ (.A1(_0887_),
    .A2(_1627_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5667_ (.A1(_1519_),
    .A2(_1632_),
    .B1(_1566_),
    .B2(_1563_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5668_ (.A1(_0745_),
    .A2(_1562_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5669_ (.A1(_1643_),
    .A2(_1644_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5670_ (.A1(_1642_),
    .A2(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5671_ (.A1(_1640_),
    .A2(_1646_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5672_ (.A1(_1560_),
    .A2(_1568_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5673_ (.A1(_1561_),
    .A2(_1567_),
    .B(_1648_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5674_ (.A1(_1631_),
    .A2(_1647_),
    .A3(_1649_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5675_ (.A1(_1626_),
    .A2(_1650_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5676_ (.I(_1651_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5677_ (.A1(_1623_),
    .A2(_1653_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5678_ (.A1(_1578_),
    .A2(_1607_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5679_ (.A1(_1575_),
    .A2(_1608_),
    .B(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5680_ (.A1(_1588_),
    .A2(_1605_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5681_ (.A1(_1584_),
    .A2(_1606_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5682_ (.A1(_1657_),
    .A2(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5683_ (.A1(_1593_),
    .A2(_1121_),
    .A3(_1592_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5684_ (.A1(_1579_),
    .A2(_1465_),
    .A3(_1595_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5685_ (.A1(_1660_),
    .A2(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5686_ (.A1(_2956_),
    .A2(_1164_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5687_ (.I(_1590_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5688_ (.I(_1476_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5689_ (.A1(_1665_),
    .A2(_1666_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5690_ (.A1(_2957_),
    .A2(_1666_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5691_ (.A1(_1591_),
    .A2(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5692_ (.A1(_1664_),
    .A2(_1667_),
    .B(_1669_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5693_ (.A1(_1593_),
    .A2(_0931_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5694_ (.A1(_1480_),
    .A2(_1664_),
    .B1(_1602_),
    .B2(_1600_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5695_ (.A1(_1599_),
    .A2(_0556_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5696_ (.A1(_1672_),
    .A2(_1673_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5697_ (.A1(_1671_),
    .A2(_1675_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5698_ (.A1(_1670_),
    .A2(_1676_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5699_ (.A1(_1596_),
    .A2(_1604_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5700_ (.A1(_1597_),
    .A2(_1603_),
    .B(_1678_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5701_ (.A1(_1662_),
    .A2(_1677_),
    .A3(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5702_ (.A1(_1659_),
    .A2(_1680_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5703_ (.I(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5704_ (.A1(_1656_),
    .A2(_1682_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5705_ (.A1(_1621_),
    .A2(_1654_),
    .A3(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5706_ (.I(_0435_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5707_ (.A1(_0392_),
    .A2(_0428_),
    .A3(_0429_),
    .B1(_0431_),
    .B2(_0357_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5708_ (.A1(_0360_),
    .A2(_0388_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5709_ (.A1(_0352_),
    .A2(_0389_),
    .A3(_0390_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5710_ (.A1(_1688_),
    .A2(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5711_ (.A1(_0371_),
    .A2(_0386_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5712_ (.A1(_0368_),
    .A2(_0387_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5713_ (.A1(_1691_),
    .A2(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5714_ (.I(_0361_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5715_ (.I(_0375_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5716_ (.A1(_1694_),
    .A2(_1695_),
    .A3(_0374_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5717_ (.A1(_0366_),
    .A2(_0363_),
    .A3(_0377_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5718_ (.A1(_1697_),
    .A2(_1698_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5719_ (.A1(_0176_),
    .A2(_0341_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5720_ (.I(_0151_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5721_ (.I(_0162_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5722_ (.A1(_1701_),
    .A2(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5723_ (.I(_0341_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5724_ (.A1(_1701_),
    .A2(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5725_ (.A1(_0373_),
    .A2(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5726_ (.A1(_1700_),
    .A2(_1703_),
    .B(_1706_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5727_ (.A1(_0365_),
    .A2(_1695_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5728_ (.A1(_0344_),
    .A2(_1700_),
    .B1(_0382_),
    .B2(_0380_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5729_ (.I(_0154_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5730_ (.A1(_0124_),
    .A2(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5731_ (.A1(_1710_),
    .A2(_1712_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5732_ (.A1(_1709_),
    .A2(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5733_ (.A1(_1708_),
    .A2(_1714_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5734_ (.A1(_0378_),
    .A2(_0385_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5735_ (.A1(_0379_),
    .A2(_0383_),
    .B(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5736_ (.A1(_1715_),
    .A2(_1717_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5737_ (.A1(_1699_),
    .A2(_1719_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5738_ (.I(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5739_ (.A1(_1693_),
    .A2(_1721_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5740_ (.A1(_1690_),
    .A2(_1722_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5741_ (.A1(_0396_),
    .A2(_0424_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5742_ (.A1(_1724_),
    .A2(_0428_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5743_ (.A1(_0408_),
    .A2(_0422_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5744_ (.A1(_0405_),
    .A2(_0423_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5745_ (.A1(_1726_),
    .A2(_1727_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5746_ (.I(_0412_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5747_ (.A1(_1730_),
    .A2(_0285_),
    .A3(_0411_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5748_ (.A1(_0398_),
    .A2(_0401_),
    .A3(_0414_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5749_ (.A1(_1731_),
    .A2(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5750_ (.A1(_0303_),
    .A2(_3257_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5751_ (.I(_3240_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5752_ (.I(_0305_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5753_ (.A1(_1735_),
    .A2(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5754_ (.I(_0303_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5755_ (.A1(_1738_),
    .A2(_1736_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5756_ (.A1(_0410_),
    .A2(_1739_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5757_ (.A1(_1734_),
    .A2(_1737_),
    .B(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5758_ (.A1(_1730_),
    .A2(_0292_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5759_ (.A1(_0307_),
    .A2(_1734_),
    .B1(_0419_),
    .B2(_0417_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5760_ (.I(_3233_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5761_ (.A1(_1745_),
    .A2(_2091_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5762_ (.A1(_1744_),
    .A2(_1746_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5763_ (.A1(_1743_),
    .A2(_1747_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5764_ (.A1(_1742_),
    .A2(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5765_ (.A1(_0415_),
    .A2(_0421_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5766_ (.A1(_0416_),
    .A2(_0420_),
    .B(_1750_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5767_ (.A1(_1733_),
    .A2(_1749_),
    .A3(_1752_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5768_ (.I(_1753_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5769_ (.A1(_1728_),
    .A2(_1754_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5770_ (.A1(_1725_),
    .A2(_1755_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5771_ (.A1(_1687_),
    .A2(_1723_),
    .A3(_1756_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5772_ (.A1(_1002_),
    .A2(_1034_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5773_ (.A1(_0969_),
    .A2(_1035_),
    .B(_1758_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5774_ (.A1(_0920_),
    .A2(_1031_),
    .A3(_1032_),
    .B1(_1005_),
    .B2(_1030_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5775_ (.A1(_1010_),
    .A2(_1028_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5776_ (.A1(_1008_),
    .A2(_1029_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5777_ (.A1(_1761_),
    .A2(_1763_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5778_ (.A1(_0882_),
    .A2(_1730_),
    .A3(_1023_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5779_ (.A1(_0888_),
    .A2(_0397_),
    .A3(_1025_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5780_ (.A1(_1765_),
    .A2(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5781_ (.A1(_3237_),
    .A2(_1336_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5782_ (.A1(_1735_),
    .A2(_1633_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5783_ (.A1(_0303_),
    .A2(_1515_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5784_ (.A1(_1014_),
    .A2(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5785_ (.A1(_1768_),
    .A2(_1769_),
    .B(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5786_ (.A1(_0412_),
    .A2(_0886_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5787_ (.A1(_0907_),
    .A2(_1768_),
    .B1(_1018_),
    .B2(_1013_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5788_ (.A1(_1745_),
    .A2(_1325_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5789_ (.A1(_1775_),
    .A2(_1776_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5790_ (.A1(_1774_),
    .A2(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5791_ (.A1(_1772_),
    .A2(_1778_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5792_ (.A1(_1020_),
    .A2(_1027_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5793_ (.A1(_1011_),
    .A2(_1019_),
    .B(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5794_ (.A1(_1767_),
    .A2(_1779_),
    .A3(_1781_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5795_ (.I(_1782_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5796_ (.A1(_1764_),
    .A2(_1783_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5797_ (.A1(_1760_),
    .A2(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5798_ (.I(_0998_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5799_ (.A1(_0972_),
    .A2(_1787_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5800_ (.A1(_0962_),
    .A2(_0999_),
    .A3(_1000_),
    .B(_1788_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5801_ (.A1(_0979_),
    .A2(_0996_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5802_ (.A1(_0976_),
    .A2(_0997_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5803_ (.A1(_1790_),
    .A2(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5804_ (.A1(_1121_),
    .A2(_1695_),
    .A3(_0983_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5805_ (.A1(_1465_),
    .A2(_0363_),
    .A3(_0985_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5806_ (.A1(_1793_),
    .A2(_1794_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5807_ (.A1(_1164_),
    .A2(_0341_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5808_ (.A1(_1666_),
    .A2(_1702_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5809_ (.A1(_1476_),
    .A2(_1704_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5810_ (.A1(_0981_),
    .A2(_1799_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5811_ (.A1(_1797_),
    .A2(_1798_),
    .B(_1800_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5812_ (.A1(_0931_),
    .A2(_0375_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5813_ (.A1(_0951_),
    .A2(_1797_),
    .B1(_0992_),
    .B2(_0989_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5814_ (.A1(_0555_),
    .A2(_1711_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5815_ (.A1(_1803_),
    .A2(_1804_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5816_ (.A1(_1802_),
    .A2(_1805_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5817_ (.A1(_1801_),
    .A2(_1807_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5818_ (.A1(_0986_),
    .A2(_0995_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5819_ (.A1(_0987_),
    .A2(_0994_),
    .B(_1809_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5820_ (.A1(_1808_),
    .A2(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5821_ (.A1(_1796_),
    .A2(_1811_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5822_ (.A1(_1789_),
    .A2(_1792_),
    .A3(_1812_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5823_ (.A1(_1786_),
    .A2(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5824_ (.A1(_1786_),
    .A2(_1813_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5825_ (.A1(_1814_),
    .A2(_1815_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5826_ (.I(_0438_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5827_ (.I(_1818_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5828_ (.A1(_1759_),
    .A2(_1816_),
    .B(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5829_ (.A1(_1759_),
    .A2(_1816_),
    .B(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5830_ (.A1(_1686_),
    .A2(_1757_),
    .B(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5831_ (.I(_3117_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5832_ (.A1(_3086_),
    .A2(_1823_),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5833_ (.A1(_3084_),
    .A2(_1824_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5834_ (.A1(_1825_),
    .A2(_3124_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5835_ (.A1(_3088_),
    .A2(_3116_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5836_ (.A1(_3086_),
    .A2(_1823_),
    .B(_1827_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5837_ (.A1(_3096_),
    .A2(_3114_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5838_ (.A1(_3094_),
    .A2(_3115_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5839_ (.A1(_2704_),
    .A2(_1627_),
    .A3(_3109_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5840_ (.A1(_0401_),
    .A2(_1546_),
    .A3(_3112_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5841_ (.A1(_1832_),
    .A2(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5842_ (.A1(_1316_),
    .A2(_3257_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5843_ (.A1(_1634_),
    .A2(_1736_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5844_ (.A1(_1513_),
    .A2(_0305_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5845_ (.A1(_3102_),
    .A2(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5846_ (.A1(_1835_),
    .A2(_1836_),
    .B(_1838_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5847_ (.A1(_1516_),
    .A2(_2708_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5848_ (.A1(_2727_),
    .A2(_1835_),
    .B1(_3104_),
    .B2(_3101_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5849_ (.A1(_3100_),
    .A2(_2080_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5850_ (.A1(_1842_),
    .A2(_1843_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5851_ (.A1(_1841_),
    .A2(_1844_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5852_ (.A1(_1840_),
    .A2(_1845_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5853_ (.A1(_3106_),
    .A2(_3113_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5854_ (.A1(_3097_),
    .A2(_3105_),
    .B(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5855_ (.A1(_1834_),
    .A2(_1846_),
    .A3(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5856_ (.A1(_1830_),
    .A2(_1831_),
    .B(_1849_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5857_ (.A1(_1830_),
    .A2(_1831_),
    .A3(_1849_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5858_ (.A1(_1851_),
    .A2(_1852_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5859_ (.A1(_1829_),
    .A2(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5860_ (.A1(_3077_),
    .A2(_3079_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5861_ (.A1(_2951_),
    .A2(_3081_),
    .B(_3080_),
    .C(_3082_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5862_ (.A1(_1855_),
    .A2(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5863_ (.A1(_3073_),
    .A2(_3076_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5864_ (.A1(_3063_),
    .A2(_3068_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5865_ (.A1(_3060_),
    .A2(_3069_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5866_ (.A1(_1859_),
    .A2(_1860_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5867_ (.A1(_3064_),
    .A2(_3067_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5868_ (.A1(_3065_),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5869_ (.A1(_3319_),
    .A2(_2863_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5870_ (.A1(_2936_),
    .A2(_2853_),
    .A3(_2810_),
    .A4(_2835_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5871_ (.A1(_0105_),
    .A2(_2811_),
    .B1(_2835_),
    .B2(_3322_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5872_ (.A1(_1866_),
    .A2(_1867_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5873_ (.A1(_1865_),
    .A2(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5874_ (.A1(_1864_),
    .A2(_1869_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5875_ (.A1(_3057_),
    .A2(_1870_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5876_ (.A1(_1862_),
    .A2(_1871_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5877_ (.A1(_3058_),
    .A2(_1873_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5878_ (.A1(_3055_),
    .A2(_3070_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5879_ (.A1(_3052_),
    .A2(_3072_),
    .B(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5880_ (.A1(_1874_),
    .A2(_1876_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5881_ (.A1(_1858_),
    .A2(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5882_ (.A1(_1857_),
    .A2(_1878_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5883_ (.A1(_1826_),
    .A2(_1854_),
    .A3(_1879_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5884_ (.A1(_0433_),
    .A2(_1880_),
    .B(_0434_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5885_ (.I(net1),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5886_ (.I(_1882_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5887_ (.A1(_1822_),
    .A2(_1881_),
    .B(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5888_ (.A1(_1617_),
    .A2(_1684_),
    .B(_1885_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5889_ (.A1(_1041_),
    .A2(_0434_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5890_ (.I(_1886_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5891_ (.A1(_1854_),
    .A2(_1879_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5892_ (.A1(_1874_),
    .A2(_1876_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5893_ (.A1(_1858_),
    .A2(_1877_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5894_ (.A1(_1857_),
    .A2(_1878_),
    .B(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5895_ (.A1(_1865_),
    .A2(_1868_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5896_ (.A1(_0329_),
    .A2(_1599_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5897_ (.A1(_0124_),
    .A2(_1590_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5898_ (.A1(_1701_),
    .A2(_2957_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5899_ (.A1(_1894_),
    .A2(_1895_),
    .A3(_1896_),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5900_ (.I(_1897_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5901_ (.A1(_1866_),
    .A2(_1892_),
    .B(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5902_ (.A1(_1866_),
    .A2(_1892_),
    .A3(_1898_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5903_ (.A1(_1899_),
    .A2(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5904_ (.I(_2957_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5905_ (.A1(_0176_),
    .A2(_1902_),
    .A3(_1870_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5906_ (.A1(_1864_),
    .A2(_1869_),
    .B(_1903_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5907_ (.A1(_1901_),
    .A2(_1905_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5908_ (.A1(_1859_),
    .A2(_1860_),
    .B(_1871_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5909_ (.A1(_3058_),
    .A2(_1873_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5910_ (.A1(_1907_),
    .A2(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5911_ (.A1(_1906_),
    .A2(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5912_ (.A1(_1889_),
    .A2(_1891_),
    .A3(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5913_ (.A1(_1829_),
    .A2(_1853_),
    .B(_1851_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5914_ (.A1(_1846_),
    .A2(_1848_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5915_ (.A1(_1846_),
    .A2(_1848_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5916_ (.A1(_1834_),
    .A2(_1913_),
    .B(_1914_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5917_ (.I(_1562_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5918_ (.A1(_1917_),
    .A2(_0399_),
    .A3(_1842_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5919_ (.A1(_1841_),
    .A2(_1844_),
    .B(_1918_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5920_ (.I(_1845_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5921_ (.A1(_1840_),
    .A2(_1920_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5922_ (.A1(_1634_),
    .A2(_2479_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5923_ (.I0(_1922_),
    .I1(_2091_),
    .S(_1838_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5924_ (.A1(_1562_),
    .A2(_0292_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5925_ (.A1(_1923_),
    .A2(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5926_ (.A1(_1837_),
    .A2(_1925_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5927_ (.A1(_1921_),
    .A2(_1927_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5928_ (.A1(_1919_),
    .A2(_1928_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5929_ (.A1(_1916_),
    .A2(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5930_ (.A1(_1916_),
    .A2(_1929_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5931_ (.A1(_1930_),
    .A2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5932_ (.A1(_1911_),
    .A2(_1912_),
    .A3(_1932_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5933_ (.A1(_1854_),
    .A2(_1879_),
    .B(_1825_),
    .C(_3124_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5934_ (.A1(_1888_),
    .A2(_1933_),
    .A3(_1934_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5935_ (.A1(_1888_),
    .A2(_1934_),
    .B(_1933_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5936_ (.A1(_1887_),
    .A2(_1935_),
    .A3(_1936_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5937_ (.A1(_0969_),
    .A2(_1035_),
    .B(_1814_),
    .C(_1758_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5938_ (.I(_1792_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5939_ (.A1(_1940_),
    .A2(_1812_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5940_ (.A1(_1940_),
    .A2(_1812_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5941_ (.A1(_1789_),
    .A2(_1941_),
    .B(_1942_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5942_ (.A1(_1796_),
    .A2(_1811_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5943_ (.A1(_1808_),
    .A2(_1810_),
    .B(_1944_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5944_ (.I(_1580_),
    .Z(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5945_ (.I(_1711_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5946_ (.A1(_1946_),
    .A2(_1947_),
    .A3(_1803_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5947_ (.A1(_1802_),
    .A2(_1805_),
    .B(_1949_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5948_ (.I(_1807_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5949_ (.A1(_1801_),
    .A2(_1951_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5950_ (.A1(_0557_),
    .A2(_1702_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5951_ (.A1(_0981_),
    .A2(_1799_),
    .B(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5952_ (.A1(_0973_),
    .A2(_1800_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5953_ (.A1(_1954_),
    .A2(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5954_ (.A1(_0932_),
    .A2(_1947_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5955_ (.A1(_1956_),
    .A2(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5956_ (.A1(_1799_),
    .A2(_1958_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5957_ (.A1(_1952_),
    .A2(_1960_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5958_ (.A1(_1950_),
    .A2(_1961_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5959_ (.A1(_1943_),
    .A2(_1945_),
    .A3(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5960_ (.A1(_1764_),
    .A2(_1783_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5961_ (.I(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5962_ (.A1(_1760_),
    .A2(_1785_),
    .B(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5963_ (.A1(_1779_),
    .A2(_1781_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5964_ (.A1(_1779_),
    .A2(_1781_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5965_ (.A1(_1767_),
    .A2(_1967_),
    .B(_1968_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5966_ (.I(_1745_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5967_ (.A1(_1971_),
    .A2(_1545_),
    .A3(_1775_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5968_ (.A1(_1774_),
    .A2(_1777_),
    .B(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5969_ (.I(_1778_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5970_ (.A1(_1772_),
    .A2(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5971_ (.A1(_3240_),
    .A2(_0745_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5972_ (.I0(_1976_),
    .I1(_0746_),
    .S(_1771_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5973_ (.A1(_1745_),
    .A2(_0887_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5974_ (.A1(_1977_),
    .A2(_1978_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5975_ (.A1(_1770_),
    .A2(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5976_ (.A1(_1975_),
    .A2(_1980_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5977_ (.A1(_1973_),
    .A2(_1982_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5978_ (.A1(_1969_),
    .A2(_1983_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5979_ (.A1(_1966_),
    .A2(_1984_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5980_ (.A1(_1963_),
    .A2(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5981_ (.A1(_1815_),
    .A2(_1939_),
    .B(_1986_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5982_ (.A1(_1815_),
    .A2(_1986_),
    .A3(_1939_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5983_ (.A1(_1819_),
    .A2(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5984_ (.A1(_1723_),
    .A2(_1756_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5985_ (.A1(_1723_),
    .A2(_1756_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5986_ (.A1(_1687_),
    .A2(_1990_),
    .B(_1991_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5987_ (.A1(_1728_),
    .A2(_1754_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5988_ (.A1(_1724_),
    .A2(_0428_),
    .B(_1755_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5989_ (.A1(_1749_),
    .A2(_1752_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5990_ (.A1(_1749_),
    .A2(_1752_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5991_ (.A1(_1733_),
    .A2(_1996_),
    .B(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5992_ (.I(_0399_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5993_ (.A1(_1971_),
    .A2(_1999_),
    .A3(_1744_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5994_ (.A1(_1743_),
    .A2(_1747_),
    .B(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5995_ (.I(_1748_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5996_ (.A1(_1742_),
    .A2(_2002_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5997_ (.A1(_3240_),
    .A2(_2091_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5998_ (.A1(_0410_),
    .A2(_1739_),
    .B(_2005_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5999_ (.A1(_2489_),
    .A2(_1741_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6000_ (.A1(_2006_),
    .A2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6001_ (.A1(_1971_),
    .A2(_2709_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6002_ (.A1(_2008_),
    .A2(_2009_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6003_ (.A1(_1739_),
    .A2(_2010_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6004_ (.A1(_2004_),
    .A2(_2011_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6005_ (.A1(_2001_),
    .A2(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6006_ (.A1(_1998_),
    .A2(_2013_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6007_ (.A1(_1994_),
    .A2(_1995_),
    .B(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6008_ (.A1(_1994_),
    .A2(_1995_),
    .A3(_2015_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6009_ (.A1(_2016_),
    .A2(_2017_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6010_ (.A1(_1693_),
    .A2(_1721_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6011_ (.A1(_1688_),
    .A2(_1689_),
    .B(_1722_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6012_ (.A1(_2019_),
    .A2(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6013_ (.I(_1719_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6014_ (.A1(_1715_),
    .A2(_1717_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6015_ (.A1(_1699_),
    .A2(_2022_),
    .B(_2023_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6016_ (.A1(_1694_),
    .A2(_1947_),
    .A3(_1710_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6017_ (.A1(_1709_),
    .A2(_1713_),
    .B(_2026_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6018_ (.I(_1714_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6019_ (.A1(_1708_),
    .A2(_2028_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6020_ (.A1(_0124_),
    .A2(_0162_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6021_ (.A1(_0373_),
    .A2(_1705_),
    .B(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6022_ (.A1(_0125_),
    .A2(_1706_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6023_ (.A1(_2031_),
    .A2(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6024_ (.A1(_0365_),
    .A2(_1711_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6025_ (.A1(_2033_),
    .A2(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6026_ (.A1(_1705_),
    .A2(_2035_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6027_ (.A1(_2029_),
    .A2(_2037_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6028_ (.A1(_2027_),
    .A2(_2038_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6029_ (.A1(_2024_),
    .A2(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6030_ (.A1(_2021_),
    .A2(_2040_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6031_ (.A1(_2018_),
    .A2(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6032_ (.A1(_1993_),
    .A2(_2042_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6033_ (.A1(_1993_),
    .A2(_2042_),
    .B(_0436_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6034_ (.A1(_1987_),
    .A2(_1989_),
    .B1(_2043_),
    .B2(_2044_),
    .C(_1039_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6035_ (.A1(_1654_),
    .A2(_1683_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6036_ (.A1(_1654_),
    .A2(_1683_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6037_ (.A1(_1621_),
    .A2(_2046_),
    .B(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6038_ (.A1(_1657_),
    .A2(_1658_),
    .B(_1680_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6039_ (.A1(_1656_),
    .A2(_1682_),
    .B(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6040_ (.A1(_1677_),
    .A2(_1679_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6041_ (.A1(_1677_),
    .A2(_1679_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6042_ (.A1(_1662_),
    .A2(_2052_),
    .B(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6043_ (.I(_1599_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6044_ (.A1(_2055_),
    .A2(_1946_),
    .A3(_1672_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6045_ (.A1(_1671_),
    .A2(_1675_),
    .B(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6046_ (.I(_1676_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6047_ (.A1(_1670_),
    .A2(_2059_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6048_ (.A1(_1590_),
    .A2(_0557_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6049_ (.A1(_1591_),
    .A2(_1668_),
    .B(_2061_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6050_ (.A1(_0973_),
    .A2(_1669_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6051_ (.A1(_2062_),
    .A2(_2063_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6052_ (.A1(_2055_),
    .A2(_0932_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6053_ (.A1(_2064_),
    .A2(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6054_ (.A1(_1668_),
    .A2(_2066_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6055_ (.A1(_2060_),
    .A2(_2067_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6056_ (.A1(_2057_),
    .A2(_2068_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6057_ (.A1(_2054_),
    .A2(_2070_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6058_ (.A1(_2054_),
    .A2(_2070_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6059_ (.A1(_2071_),
    .A2(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6060_ (.A1(_2051_),
    .A2(_2073_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6061_ (.A1(_1624_),
    .A2(_1625_),
    .B(_1650_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6062_ (.A1(_1623_),
    .A2(_1653_),
    .B(_2075_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6063_ (.A1(_1647_),
    .A2(_1649_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6064_ (.A1(_1647_),
    .A2(_1649_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6065_ (.A1(_1631_),
    .A2(_2077_),
    .B(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6066_ (.I(_1545_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6067_ (.A1(_2081_),
    .A2(_1917_),
    .A3(_1643_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6068_ (.A1(_1642_),
    .A2(_1645_),
    .B(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6069_ (.I(_1646_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6070_ (.A1(_1640_),
    .A2(_2084_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6071_ (.A1(_0746_),
    .A2(_1634_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6072_ (.A1(_1556_),
    .A2(_1638_),
    .B(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6073_ (.A1(_0882_),
    .A2(_1639_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6074_ (.A1(_2087_),
    .A2(_2088_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6075_ (.A1(_0888_),
    .A2(_1917_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6076_ (.A1(_2089_),
    .A2(_2090_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6077_ (.A1(_1638_),
    .A2(_2092_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6078_ (.A1(_2085_),
    .A2(_2093_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6079_ (.A1(_2083_),
    .A2(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6080_ (.A1(_2079_),
    .A2(_2095_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6081_ (.A1(_2079_),
    .A2(_2095_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6082_ (.A1(_2096_),
    .A2(_2097_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6083_ (.A1(_2076_),
    .A2(_2098_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6084_ (.A1(_2049_),
    .A2(_2074_),
    .A3(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6085_ (.A1(_1043_),
    .A2(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6086_ (.A1(_1938_),
    .A2(_2045_),
    .B(_2101_),
    .C(_1614_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6087_ (.A1(_1912_),
    .A2(_1932_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6088_ (.A1(_1912_),
    .A2(_1932_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6089_ (.A1(_1911_),
    .A2(_2103_),
    .A3(_2104_),
    .B(_1935_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6090_ (.A1(_1889_),
    .A2(_1910_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6091_ (.A1(_1889_),
    .A2(_1910_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6092_ (.A1(_1891_),
    .A2(_2106_),
    .B(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6093_ (.A1(_1906_),
    .A2(_1909_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6094_ (.I(_1901_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6095_ (.A1(_2110_),
    .A2(_1905_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6096_ (.A1(_1899_),
    .A2(_2111_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6097_ (.A1(_1694_),
    .A2(_2055_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6098_ (.A1(_0365_),
    .A2(_1665_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6099_ (.A1(_1894_),
    .A2(_1895_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6100_ (.A1(_2114_),
    .A2(_2115_),
    .B1(_1896_),
    .B2(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6101_ (.A1(_0361_),
    .A2(_1902_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6102_ (.A1(_2115_),
    .A2(_2118_),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6103_ (.A1(_2117_),
    .A2(_2119_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6104_ (.A1(_2113_),
    .A2(_2120_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6105_ (.A1(_2109_),
    .A2(_2121_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6106_ (.A1(_2108_),
    .A2(_2122_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6107_ (.A1(_1912_),
    .A2(_1932_),
    .B(_1930_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6108_ (.A1(_1921_),
    .A2(_1927_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6109_ (.A1(_1919_),
    .A2(_1928_),
    .B(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6110_ (.A1(_1999_),
    .A2(_1838_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6111_ (.A1(_1923_),
    .A2(_1924_),
    .B(_2128_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6112_ (.A1(_1837_),
    .A2(_1925_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6113_ (.A1(_1637_),
    .A2(_0285_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6114_ (.A1(_1635_),
    .A2(_0401_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6115_ (.A1(_2131_),
    .A2(_2132_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6116_ (.A1(_2130_),
    .A2(_2133_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6117_ (.A1(_2129_),
    .A2(_2135_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6118_ (.A1(_2127_),
    .A2(_2136_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6119_ (.A1(_2125_),
    .A2(_2137_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6120_ (.A1(_2124_),
    .A2(_2138_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6121_ (.A1(_2105_),
    .A2(_2139_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6122_ (.A1(_2105_),
    .A2(_2139_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6123_ (.A1(_1887_),
    .A2(_2140_),
    .A3(_2141_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6124_ (.A1(_1963_),
    .A2(_1985_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6125_ (.A1(_1945_),
    .A2(_1962_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6126_ (.A1(_1945_),
    .A2(_1962_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6127_ (.A1(_1943_),
    .A2(_2144_),
    .B(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6128_ (.A1(_1952_),
    .A2(_1960_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6129_ (.A1(_1950_),
    .A2(_1961_),
    .B(_2148_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6130_ (.A1(_1956_),
    .A2(_1957_),
    .B(_1955_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6131_ (.A1(_1799_),
    .A2(_1958_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6132_ (.I(_1704_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6133_ (.I(_1702_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6134_ (.A1(_1580_),
    .A2(_2152_),
    .B1(_2153_),
    .B2(_1465_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6135_ (.A1(_1124_),
    .A2(_2152_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6136_ (.A1(_1953_),
    .A2(_2155_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6137_ (.A1(_2154_),
    .A2(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6138_ (.A1(_2151_),
    .A2(_2158_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6139_ (.A1(_2150_),
    .A2(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6140_ (.A1(_2149_),
    .A2(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6141_ (.A1(_2147_),
    .A2(_2161_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6142_ (.I(_1969_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6143_ (.A1(_2163_),
    .A2(_1983_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6144_ (.A1(_1966_),
    .A2(_1984_),
    .B(_2164_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6145_ (.A1(_1975_),
    .A2(_1980_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6146_ (.A1(_1973_),
    .A2(_1982_),
    .B(_2166_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6147_ (.A1(_2081_),
    .A2(_1771_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6148_ (.A1(_1977_),
    .A2(_1978_),
    .B(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6149_ (.A1(_1770_),
    .A2(_1979_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6150_ (.I(_1738_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6151_ (.I(_1735_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6152_ (.A1(_2172_),
    .A2(_1292_),
    .B1(_1294_),
    .B2(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6153_ (.A1(_1738_),
    .A2(_0889_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6154_ (.A1(_1976_),
    .A2(_2175_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6155_ (.A1(_2174_),
    .A2(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6156_ (.A1(_2171_),
    .A2(_2177_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6157_ (.A1(_2170_),
    .A2(_2179_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6158_ (.A1(_2168_),
    .A2(_2180_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6159_ (.A1(_2165_),
    .A2(_2181_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6160_ (.A1(_2162_),
    .A2(_2182_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6161_ (.A1(_2143_),
    .A2(_1988_),
    .B(_2183_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6162_ (.I(_1818_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6163_ (.A1(_2143_),
    .A2(_1988_),
    .A3(_2183_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6164_ (.A1(_2185_),
    .A2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6165_ (.A1(_2018_),
    .A2(_2041_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6166_ (.A1(_1993_),
    .A2(_2042_),
    .B(_2188_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6167_ (.A1(_1998_),
    .A2(_2013_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6168_ (.A1(_2004_),
    .A2(_2011_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6169_ (.A1(_2001_),
    .A2(_2012_),
    .B(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6170_ (.A1(_2008_),
    .A2(_2009_),
    .B(_2007_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6171_ (.A1(_1739_),
    .A2(_2010_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6172_ (.A1(_2172_),
    .A2(_1999_),
    .B1(_0402_),
    .B2(_2173_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6173_ (.A1(_1738_),
    .A2(_1735_),
    .A3(_0399_),
    .A4(_0402_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6174_ (.A1(_2196_),
    .A2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6175_ (.A1(_2195_),
    .A2(_2198_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6176_ (.A1(_2194_),
    .A2(_2199_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6177_ (.A1(_2193_),
    .A2(_2201_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6178_ (.A1(_2191_),
    .A2(_2016_),
    .B(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6179_ (.A1(_2191_),
    .A2(_2016_),
    .A3(_2202_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6180_ (.A1(_2203_),
    .A2(_2204_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6181_ (.A1(_2024_),
    .A2(_2039_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6182_ (.A1(_2019_),
    .A2(_2020_),
    .B(_2040_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6183_ (.A1(_2029_),
    .A2(_2037_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6184_ (.A1(_2027_),
    .A2(_2038_),
    .B(_2208_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6185_ (.A1(_2033_),
    .A2(_2034_),
    .B(_2032_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6186_ (.A1(_1705_),
    .A2(_2035_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6187_ (.A1(_0361_),
    .A2(_1704_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6188_ (.A1(_0366_),
    .A2(_2153_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6189_ (.A1(_2213_),
    .A2(_2214_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6190_ (.A1(_2212_),
    .A2(_2215_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6191_ (.A1(_2210_),
    .A2(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6192_ (.A1(_2209_),
    .A2(_2217_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6193_ (.A1(_2206_),
    .A2(_2207_),
    .B(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6194_ (.A1(_2206_),
    .A2(_2207_),
    .A3(_2218_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6195_ (.A1(_2219_),
    .A2(_2220_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6196_ (.A1(_2205_),
    .A2(_2221_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6197_ (.A1(_2190_),
    .A2(_2223_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6198_ (.A1(_2190_),
    .A2(_2223_),
    .B(_1686_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6199_ (.I(_1615_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6200_ (.A1(_2184_),
    .A2(_2187_),
    .B1(_2224_),
    .B2(_2225_),
    .C(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6201_ (.A1(_2074_),
    .A2(_2099_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6202_ (.A1(_2074_),
    .A2(_2099_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6203_ (.A1(_2049_),
    .A2(_2228_),
    .B(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6204_ (.A1(_2051_),
    .A2(_2073_),
    .B(_2071_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6205_ (.A1(_2060_),
    .A2(_2067_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6206_ (.A1(_2057_),
    .A2(_2068_),
    .B(_2232_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6207_ (.A1(_2064_),
    .A2(_2065_),
    .B(_2063_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6208_ (.A1(_1668_),
    .A2(_2066_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6209_ (.A1(_1902_),
    .A2(_1580_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6210_ (.A1(_1665_),
    .A2(_1582_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6211_ (.A1(_2237_),
    .A2(_2238_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6212_ (.A1(_2236_),
    .A2(_2239_),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6213_ (.A1(_2235_),
    .A2(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6214_ (.A1(_2234_),
    .A2(_2241_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6215_ (.A1(_2231_),
    .A2(_2242_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6216_ (.A1(_2076_),
    .A2(_2098_),
    .B(_2096_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6217_ (.A1(_2085_),
    .A2(_2093_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6218_ (.A1(_2083_),
    .A2(_2094_),
    .B(_2246_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6219_ (.A1(_2089_),
    .A2(_2090_),
    .B(_2088_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6220_ (.A1(_1638_),
    .A2(_2092_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6221_ (.A1(_1545_),
    .A2(_1637_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6222_ (.A1(_1548_),
    .A2(_1635_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6223_ (.A1(_2250_),
    .A2(_2251_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6224_ (.A1(_2249_),
    .A2(_2252_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6225_ (.A1(_2248_),
    .A2(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6226_ (.A1(_2247_),
    .A2(_2254_),
    .Z(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6227_ (.A1(_2245_),
    .A2(_2256_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6228_ (.A1(_2243_),
    .A2(_2257_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6229_ (.A1(_2230_),
    .A2(_2258_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6230_ (.A1(_1043_),
    .A2(_2259_),
    .B(_1884_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6231_ (.A1(_2142_),
    .A2(_2227_),
    .B(_2260_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6232_ (.I(_1882_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6233_ (.A1(_2205_),
    .A2(_2221_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6234_ (.A1(_2190_),
    .A2(_2223_),
    .B(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6235_ (.A1(_2193_),
    .A2(_2201_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6236_ (.A1(_2195_),
    .A2(_2198_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6237_ (.A1(_2194_),
    .A2(_2199_),
    .B(_2266_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6238_ (.I(_0402_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6239_ (.A1(_2172_),
    .A2(_2268_),
    .A3(_2005_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6240_ (.A1(_2267_),
    .A2(_2269_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6241_ (.A1(_2264_),
    .A2(_2203_),
    .B(_2270_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6242_ (.A1(_2264_),
    .A2(_2203_),
    .A3(_2270_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6243_ (.A1(_2271_),
    .A2(_2272_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6244_ (.A1(_2212_),
    .A2(_2215_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6245_ (.A1(_2210_),
    .A2(_2216_),
    .B(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6246_ (.I(_0366_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6247_ (.A1(_2277_),
    .A2(_2152_),
    .A3(_2030_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6248_ (.A1(_2275_),
    .A2(_2278_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6249_ (.A1(_2209_),
    .A2(_2217_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6250_ (.A1(_2280_),
    .A2(_2219_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6251_ (.A1(_2279_),
    .A2(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6252_ (.A1(_2273_),
    .A2(_2282_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6253_ (.A1(_2263_),
    .A2(_2283_),
    .B(_0436_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6254_ (.A1(_2263_),
    .A2(_2283_),
    .B(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6255_ (.A1(_2162_),
    .A2(_2182_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6256_ (.A1(_2286_),
    .A2(_2184_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6257_ (.A1(_2151_),
    .A2(_2158_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6258_ (.A1(_2150_),
    .A2(_2159_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6259_ (.A1(_2289_),
    .A2(_2290_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6260_ (.A1(_1946_),
    .A2(_2153_),
    .B(_2155_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6261_ (.A1(_2291_),
    .A2(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6262_ (.A1(_2149_),
    .A2(_2160_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6263_ (.A1(_2147_),
    .A2(_2161_),
    .B(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6264_ (.A1(_2293_),
    .A2(_2295_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6265_ (.A1(_2171_),
    .A2(_2177_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6266_ (.A1(_2170_),
    .A2(_2179_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6267_ (.A1(_2297_),
    .A2(_2299_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6268_ (.A1(_2173_),
    .A2(_2081_),
    .B(_2175_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6269_ (.A1(_2300_),
    .A2(_2301_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6270_ (.A1(_2168_),
    .A2(_2180_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6271_ (.A1(_2165_),
    .A2(_2181_),
    .B(_2303_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6272_ (.A1(_2302_),
    .A2(_2304_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6273_ (.A1(_2296_),
    .A2(_2305_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6274_ (.A1(_2288_),
    .A2(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6275_ (.A1(_2124_),
    .A2(_2138_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6276_ (.A1(_2105_),
    .A2(_2139_),
    .B(_2308_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6277_ (.A1(_1906_),
    .A2(_1909_),
    .A3(_2121_),
    .B1(_2122_),
    .B2(_2108_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6278_ (.A1(_2111_),
    .A2(_2120_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6279_ (.I(_1902_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6280_ (.A1(_2277_),
    .A2(_2313_),
    .A3(_1895_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6281_ (.A1(_2117_),
    .A2(_2119_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6282_ (.A1(_1899_),
    .A2(_2120_),
    .B(_2315_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6283_ (.A1(_2314_),
    .A2(_2316_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6284_ (.A1(_2312_),
    .A2(_2317_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6285_ (.A1(_2311_),
    .A2(_2318_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6286_ (.A1(_2130_),
    .A2(_2133_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6287_ (.A1(_2129_),
    .A2(_2135_),
    .B(_2321_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6288_ (.I(_1637_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6289_ (.A1(_2323_),
    .A2(_2268_),
    .A3(_1922_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6290_ (.A1(_2322_),
    .A2(_2324_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6291_ (.I(_2325_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6292_ (.A1(_2127_),
    .A2(_2136_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6293_ (.A1(_2125_),
    .A2(_2137_),
    .B(_2327_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6294_ (.A1(_2326_),
    .A2(_2328_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6295_ (.A1(_2310_),
    .A2(_2319_),
    .A3(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6296_ (.A1(_0440_),
    .A2(_2307_),
    .B1(_2330_),
    .B2(_1887_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6297_ (.A1(_1043_),
    .A2(_2285_),
    .A3(_2332_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6298_ (.A1(_2236_),
    .A2(_2239_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6299_ (.A1(_2235_),
    .A2(_2240_),
    .B(_2334_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6300_ (.A1(_2313_),
    .A2(_1582_),
    .A3(_2061_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6301_ (.A1(_2335_),
    .A2(_2336_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6302_ (.A1(_2234_),
    .A2(_2241_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6303_ (.A1(_2231_),
    .A2(_2242_),
    .B(_2338_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6304_ (.A1(_2337_),
    .A2(_2339_),
    .Z(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6305_ (.A1(_2249_),
    .A2(_2252_),
    .Z(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6306_ (.A1(_2248_),
    .A2(_2253_),
    .B(_2341_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6307_ (.A1(_1548_),
    .A2(_2323_),
    .A3(_2086_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6308_ (.A1(_2343_),
    .A2(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6309_ (.A1(_2247_),
    .A2(_2254_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6310_ (.A1(_2245_),
    .A2(_2256_),
    .B(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6311_ (.A1(_2345_),
    .A2(_2347_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6312_ (.A1(_2340_),
    .A2(_2348_),
    .Z(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6313_ (.A1(_2243_),
    .A2(_2257_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6314_ (.A1(_2230_),
    .A2(_2258_),
    .B(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6315_ (.A1(_2349_),
    .A2(_2351_),
    .B(_1042_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6316_ (.A1(_2349_),
    .A2(_2351_),
    .B(_2352_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6317_ (.A1(_2261_),
    .A2(_2333_),
    .A3(_2354_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6318_ (.I(_2355_),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6319_ (.A1(_2319_),
    .A2(_2329_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6320_ (.A1(_2319_),
    .A2(_2329_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6321_ (.A1(_2310_),
    .A2(_2356_),
    .B(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6322_ (.I(_2316_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6323_ (.A1(_2277_),
    .A2(_2313_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6324_ (.A1(_1895_),
    .A2(_2359_),
    .B(_2360_),
    .ZN(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6325_ (.A1(_2312_),
    .A2(_2317_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6326_ (.A1(_2311_),
    .A2(_2318_),
    .B(_2361_),
    .C(_2362_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6327_ (.A1(_2326_),
    .A2(_2328_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6328_ (.A1(_2323_),
    .A2(_2268_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6329_ (.A1(_1922_),
    .A2(_2322_),
    .B(_2366_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6330_ (.A1(_2365_),
    .A2(_2367_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6331_ (.A1(_2364_),
    .A2(_2368_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6332_ (.A1(_2358_),
    .A2(_2369_),
    .B(_3123_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6333_ (.A1(_2358_),
    .A2(_2369_),
    .B(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6334_ (.A1(_2273_),
    .A2(_2282_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6335_ (.A1(_2263_),
    .A2(_2283_),
    .B(_2372_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6336_ (.A1(_2267_),
    .A2(_2269_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6337_ (.A1(_2197_),
    .A2(_2375_),
    .A3(_2271_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6338_ (.A1(_2280_),
    .A2(_2219_),
    .B(_2279_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6339_ (.A1(_2213_),
    .A2(_2214_),
    .B1(_2275_),
    .B2(_2278_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6340_ (.A1(_2377_),
    .A2(_2378_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6341_ (.A1(_2376_),
    .A2(_2379_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6342_ (.A1(_2373_),
    .A2(_2380_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6343_ (.A1(_2373_),
    .A2(_2380_),
    .B(_1686_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6344_ (.A1(_2296_),
    .A2(_2305_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6345_ (.A1(_2286_),
    .A2(_2184_),
    .B(_2306_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6346_ (.A1(_2291_),
    .A2(_2292_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6347_ (.A1(_2293_),
    .A2(_2295_),
    .B(_2386_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6348_ (.A1(_2157_),
    .A2(_2387_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6349_ (.A1(_2300_),
    .A2(_2301_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6350_ (.A1(_2302_),
    .A2(_2304_),
    .B(_2389_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6351_ (.A1(_2176_),
    .A2(_2390_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6352_ (.A1(_2388_),
    .A2(_2391_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6353_ (.A1(_2383_),
    .A2(_2384_),
    .B(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6354_ (.A1(_2383_),
    .A2(_2384_),
    .A3(_2392_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6355_ (.A1(_2185_),
    .A2(_2394_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6356_ (.A1(_2381_),
    .A2(_2382_),
    .B1(_2393_),
    .B2(_2395_),
    .C(_2226_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6357_ (.A1(_2337_),
    .A2(_2339_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6358_ (.A1(_2237_),
    .A2(_2238_),
    .B1(_2335_),
    .B2(_2336_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6359_ (.A1(_2398_),
    .A2(_2399_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6360_ (.A1(_2345_),
    .A2(_2347_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6361_ (.A1(_2250_),
    .A2(_2251_),
    .B1(_2343_),
    .B2(_2344_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6362_ (.A1(_2401_),
    .A2(_2402_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6363_ (.A1(_2400_),
    .A2(_2403_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6364_ (.A1(_2340_),
    .A2(_2348_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6365_ (.A1(_2340_),
    .A2(_2348_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6366_ (.A1(_2405_),
    .A2(_2351_),
    .B(_2406_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6367_ (.A1(_2404_),
    .A2(_2408_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6368_ (.I(_1038_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6369_ (.A1(_2404_),
    .A2(_2408_),
    .B(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6370_ (.A1(_2409_),
    .A2(_2411_),
    .B(_1884_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6371_ (.A1(_2371_),
    .A2(_2397_),
    .B(_2412_),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6372_ (.A1(_2364_),
    .A2(_2368_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6373_ (.A1(_2388_),
    .A2(_2391_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6374_ (.A1(_1041_),
    .A2(_2393_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6375_ (.A1(_2376_),
    .A2(_2379_),
    .B(_0433_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6376_ (.A1(_2373_),
    .A2(_2380_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6377_ (.A1(_2414_),
    .A2(_2415_),
    .B1(_2416_),
    .B2(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6378_ (.A1(_2405_),
    .A2(_2351_),
    .B1(_2400_),
    .B2(_2403_),
    .C(_2406_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6379_ (.A1(_2400_),
    .A2(_2403_),
    .B(_1615_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6380_ (.I(_1882_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6381_ (.A1(_2420_),
    .A2(_2421_),
    .B(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6382_ (.A1(_2413_),
    .A2(_2370_),
    .B1(_2419_),
    .B2(_0434_),
    .C(_2423_),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6383_ (.A1(_1435_),
    .A2(_3209_),
    .B1(_0128_),
    .B2(_1434_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6384_ (.A1(_0858_),
    .A2(_0440_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6385_ (.A1(_1041_),
    .A2(_3120_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6386_ (.I(_2426_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6387_ (.A1(_3289_),
    .A2(_0208_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6388_ (.A1(_0250_),
    .A2(_2428_),
    .A3(_2429_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6389_ (.A1(_1685_),
    .A2(_2761_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6390_ (.A1(_2998_),
    .A2(_1886_),
    .A3(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6391_ (.A1(_2424_),
    .A2(_2425_),
    .B(_2430_),
    .C(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6392_ (.A1(_1126_),
    .A2(_1434_),
    .B1(_1435_),
    .B2(_1295_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6393_ (.A1(_2410_),
    .A2(_1436_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6394_ (.A1(_2434_),
    .A2(_2435_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6395_ (.A1(_2433_),
    .A2(_2436_),
    .B(_2261_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6396_ (.I(_2437_),
    .ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6397_ (.A1(_1428_),
    .A2(_1431_),
    .A3(_1436_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6398_ (.A1(_0250_),
    .A2(_0259_),
    .B(_0435_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6399_ (.A1(_0250_),
    .A2(_0259_),
    .B(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6400_ (.A1(_3007_),
    .A2(_3013_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6401_ (.A1(_2442_),
    .A2(_2999_),
    .A3(_3014_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6402_ (.A1(_2442_),
    .A2(_3014_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6403_ (.A1(_2998_),
    .A2(_2444_),
    .B(_3122_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6404_ (.A1(_0858_),
    .A2(_0859_),
    .B(_1819_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6405_ (.A1(_2443_),
    .A2(_2445_),
    .B1(_2446_),
    .B2(_0860_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6406_ (.A1(_1042_),
    .A2(_2441_),
    .A3(_2447_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6407_ (.A1(_2261_),
    .A2(_2449_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6408_ (.A1(_1617_),
    .A2(_2439_),
    .B(_2450_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6409_ (.A1(_1438_),
    .A2(_1441_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6410_ (.A1(_0261_),
    .A2(_0264_),
    .B(_2428_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6411_ (.A1(_0261_),
    .A2(_0264_),
    .B(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6412_ (.A1(_2442_),
    .A2(_2443_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6413_ (.A1(_3017_),
    .A2(_3018_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6414_ (.A1(_2454_),
    .A2(_2455_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6415_ (.A1(_2454_),
    .A2(_2455_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6416_ (.A1(_2457_),
    .A2(_1886_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6417_ (.A1(_0857_),
    .A2(_0860_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6418_ (.A1(_2460_),
    .A2(_0863_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6419_ (.A1(_2456_),
    .A2(_2459_),
    .B1(_2461_),
    .B2(_2185_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6420_ (.A1(_1616_),
    .A2(_2453_),
    .A3(_2462_),
    .B(_2422_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6421_ (.A1(_1617_),
    .A2(_2451_),
    .B(_2463_),
    .ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6422_ (.A1(_0266_),
    .A2(_0267_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6423_ (.A1(_0268_),
    .A2(_1686_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6424_ (.A1(_2464_),
    .A2(_2465_),
    .B(_2410_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6425_ (.A1(_3023_),
    .A2(_3024_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6426_ (.A1(_2467_),
    .A2(_3021_),
    .A3(_3025_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6427_ (.A1(_3020_),
    .A2(_2457_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6428_ (.A1(_2467_),
    .A2(_3025_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6429_ (.A1(_2470_),
    .A2(_2471_),
    .B(_3122_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6430_ (.A1(_0847_),
    .A2(_0864_),
    .A3(_0866_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6431_ (.A1(_1819_),
    .A2(_2473_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6432_ (.A1(_2469_),
    .A2(_2472_),
    .B1(_2474_),
    .B2(_0867_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6433_ (.A1(_1425_),
    .A2(_1443_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6434_ (.A1(_1445_),
    .A2(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6435_ (.I(_1039_),
    .Z(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6436_ (.A1(_2466_),
    .A2(_2475_),
    .B1(_2477_),
    .B2(_2478_),
    .C(_1613_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6437_ (.A1(_1424_),
    .A2(_1445_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6438_ (.A1(_2480_),
    .A2(_1446_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6439_ (.A1(_0269_),
    .A2(_0249_),
    .A3(_0268_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6440_ (.A1(_0436_),
    .A2(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6441_ (.A1(_3027_),
    .A2(_3030_),
    .B(_3121_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6442_ (.A1(_3027_),
    .A2(_3030_),
    .B(_2484_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6443_ (.A1(_0868_),
    .A2(_0841_),
    .A3(_0867_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6444_ (.A1(_0869_),
    .A2(_1818_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6445_ (.A1(_2486_),
    .A2(_2487_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6446_ (.A1(_2485_),
    .A2(_2488_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6447_ (.A1(_0270_),
    .A2(_2483_),
    .B(_2490_),
    .C(_1039_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6448_ (.A1(_2478_),
    .A2(_2481_),
    .B(_2491_),
    .C(_1614_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6449_ (.A1(_1418_),
    .A2(_1447_),
    .A3(_1448_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6450_ (.A1(_1449_),
    .A2(_2492_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6451_ (.A1(_3032_),
    .A2(_3033_),
    .B(_1886_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6452_ (.A1(_3034_),
    .A2(_2494_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6453_ (.A1(_0837_),
    .A2(_0869_),
    .A3(_0870_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6454_ (.A1(_0871_),
    .A2(_0439_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6455_ (.A1(_0271_),
    .A2(_0272_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6456_ (.A1(_0273_),
    .A2(_2428_),
    .A3(_2498_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6457_ (.A1(_2496_),
    .A2(_2497_),
    .B(_1042_),
    .C(_2500_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6458_ (.A1(_2495_),
    .A2(_2501_),
    .B(_2422_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6459_ (.A1(_1617_),
    .A2(_2493_),
    .B(_2502_),
    .ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6460_ (.A1(_2997_),
    .A2(_3034_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6461_ (.A1(_3037_),
    .A2(_3039_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6462_ (.A1(_2503_),
    .A2(_2504_),
    .B(_3123_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6463_ (.A1(_2503_),
    .A2(_2504_),
    .B(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6464_ (.I(_0874_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6465_ (.A1(_0826_),
    .A2(_2507_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6466_ (.A1(_0873_),
    .A2(_2508_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6467_ (.A1(_0236_),
    .A2(_0237_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6468_ (.A1(_0274_),
    .A2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6469_ (.A1(_0440_),
    .A2(_2510_),
    .B1(_2512_),
    .B2(_2428_),
    .C(_2226_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6470_ (.A1(_1405_),
    .A2(_1406_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6471_ (.A1(_1408_),
    .A2(_1407_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6472_ (.A1(_2514_),
    .A2(_2515_),
    .A3(_1450_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6473_ (.A1(_2226_),
    .A2(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6474_ (.A1(_1884_),
    .A2(_2517_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6475_ (.A1(_2506_),
    .A2(_2513_),
    .B(_2518_),
    .ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6476_ (.A1(_3042_),
    .A2(_3044_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6477_ (.A1(_3042_),
    .A2(_3044_),
    .B(_1887_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6478_ (.A1(_0821_),
    .A2(_0822_),
    .A3(_0875_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6479_ (.A1(_0236_),
    .A2(_0275_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6480_ (.A1(_0229_),
    .A2(_0230_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6481_ (.A1(_2523_),
    .A2(_2524_),
    .B(_2426_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6482_ (.A1(_2523_),
    .A2(_2524_),
    .B(_2525_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6483_ (.A1(_0439_),
    .A2(_2522_),
    .B(_2526_),
    .C(_1615_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6484_ (.A1(_2520_),
    .A2(_2521_),
    .B(_2527_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6485_ (.A1(_1404_),
    .A2(_1452_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6486_ (.A1(_1453_),
    .A2(_1452_),
    .B(_1454_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6487_ (.A1(_2529_),
    .A2(_2531_),
    .B(_1616_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6488_ (.A1(_2261_),
    .A2(_2528_),
    .A3(_2532_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6489_ (.I(_2533_),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6490_ (.A1(_1216_),
    .A2(_1391_),
    .A3(_1454_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6491_ (.A1(_0228_),
    .A2(_0277_),
    .B(_2426_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6492_ (.A1(_0228_),
    .A2(_0277_),
    .B(_2535_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6493_ (.A1(_3045_),
    .A2(_3046_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6494_ (.A1(_0623_),
    .A2(_0819_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6495_ (.A1(_2538_),
    .A2(_0820_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6496_ (.A1(_0823_),
    .A2(_0875_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6497_ (.A1(_0821_),
    .A2(_0822_),
    .B(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6498_ (.A1(_2539_),
    .A2(_2542_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6499_ (.A1(_0439_),
    .A2(_2543_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6500_ (.A1(_2539_),
    .A2(_2542_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6501_ (.A1(_3047_),
    .A2(_3122_),
    .A3(_2537_),
    .B1(_2544_),
    .B2(_2545_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6502_ (.A1(_2410_),
    .A2(_2536_),
    .A3(_2546_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6503_ (.A1(_2478_),
    .A2(_2534_),
    .B(_2547_),
    .C(_1614_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6504_ (.A1(_1496_),
    .A2(_1536_),
    .A3(_1457_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6505_ (.A1(_0279_),
    .A2(_0355_),
    .B(_2426_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6506_ (.A1(_0279_),
    .A2(_0355_),
    .B(_2549_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6507_ (.A1(_2990_),
    .A2(_3047_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6508_ (.A1(_2552_),
    .A2(_3048_),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6509_ (.A1(_2552_),
    .A2(_3048_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6510_ (.A1(_0879_),
    .A2(_0967_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6511_ (.A1(_2553_),
    .A2(_3123_),
    .A3(_2554_),
    .B1(_2555_),
    .B2(_2185_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6512_ (.A1(_1616_),
    .A2(_2551_),
    .A3(_2556_),
    .B(_2422_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6513_ (.A1(_2478_),
    .A2(_2548_),
    .B(_2557_),
    .ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6514_ (.I(net7),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6515_ (.I(net5),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6516_ (.A1(_1613_),
    .A2(net4),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6517_ (.A1(net6),
    .A2(_2559_),
    .A3(_2561_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6518_ (.I(_2562_),
    .Z(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6519_ (.I0(_3004_),
    .I1(_2558_),
    .S(_2563_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6520_ (.I(_2564_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6521_ (.I(net8),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6522_ (.I0(_2959_),
    .I1(_2565_),
    .S(_2563_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6523_ (.I(_2566_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6524_ (.I(net9),
    .Z(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6525_ (.I0(_2784_),
    .I1(_2567_),
    .S(_2563_),
    .Z(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6526_ (.I(_2568_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6527_ (.I(net10),
    .Z(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6528_ (.I0(_3311_),
    .I1(_2570_),
    .S(_2563_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6529_ (.I(_2571_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6530_ (.I(net11),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6531_ (.I(_2562_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6532_ (.I0(_0176_),
    .I1(_2572_),
    .S(_2573_),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6533_ (.I(_2574_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6534_ (.I(net12),
    .Z(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6535_ (.I0(_1701_),
    .I1(_2575_),
    .S(_2573_),
    .Z(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6536_ (.I(_2576_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6537_ (.I(net13),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6538_ (.I0(_1694_),
    .I1(_2578_),
    .S(_2573_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6539_ (.I(_2579_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6540_ (.I(net14),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6541_ (.I0(_2277_),
    .I1(_2580_),
    .S(_2573_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6542_ (.I(_2581_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6543_ (.A1(_1882_),
    .A2(net4),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6544_ (.A1(net6),
    .A2(_2559_),
    .A3(_2582_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6545_ (.I(_2583_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6546_ (.I0(_1434_),
    .I1(_2558_),
    .S(_2584_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6547_ (.I(_2586_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6548_ (.I0(_0848_),
    .I1(_2565_),
    .S(_2584_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6549_ (.I(_2587_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6550_ (.I0(_0946_),
    .I1(_2567_),
    .S(_2584_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6551_ (.I(_2588_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6552_ (.I0(_1045_),
    .I1(_2570_),
    .S(_2584_),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6553_ (.I(_2589_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6554_ (.I(_2583_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6555_ (.I0(_1164_),
    .I1(_2572_),
    .S(_2590_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6556_ (.I(_2591_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6557_ (.I0(_1666_),
    .I1(_2575_),
    .S(_2590_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6558_ (.I(_2593_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6559_ (.I0(_1946_),
    .I1(_2578_),
    .S(_2590_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6560_ (.I(_2594_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6561_ (.I0(_1582_),
    .I1(_2580_),
    .S(_2590_),
    .Z(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6562_ (.I(_2595_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6563_ (.I(net7),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6564_ (.I(net6),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6565_ (.A1(_2597_),
    .A2(_2559_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6566_ (.A1(_2561_),
    .A2(_2598_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6567_ (.I(_2600_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6568_ (.I0(_2596_),
    .I1(_3011_),
    .S(_2601_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6569_ (.I(_2602_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6570_ (.I(net8),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6571_ (.I0(_2603_),
    .I1(_3009_),
    .S(_2601_),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6572_ (.I(_2604_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6573_ (.I(net9),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6574_ (.I0(_2605_),
    .I1(_3247_),
    .S(_2601_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6575_ (.I(_2606_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6576_ (.I(net10),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6577_ (.I0(_2608_),
    .I1(_3128_),
    .S(_2601_),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6578_ (.I(_2609_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6579_ (.I(net11),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6580_ (.I(_2600_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6581_ (.I0(_2610_),
    .I1(_3257_),
    .S(_2611_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6582_ (.I(_2612_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6583_ (.I(net12),
    .Z(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6584_ (.I0(_2613_),
    .I1(_1736_),
    .S(_2611_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6585_ (.I(_2614_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6586_ (.I(net13),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6587_ (.I0(_2616_),
    .I1(_1999_),
    .S(_2611_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6588_ (.I(_2617_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6589_ (.I(net14),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6590_ (.I0(_2618_),
    .I1(_2268_),
    .S(_2611_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6591_ (.I(_2619_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6592_ (.A1(_2582_),
    .A2(_2598_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6593_ (.I(_2620_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6594_ (.I0(_2596_),
    .I1(_1435_),
    .S(_2621_),
    .Z(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6595_ (.I(_2622_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6596_ (.I0(_2603_),
    .I1(_0853_),
    .S(_2621_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6597_ (.I(_2624_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6598_ (.I0(_2605_),
    .I1(_0909_),
    .S(_2621_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6599_ (.I(_2625_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6600_ (.I0(_2608_),
    .I1(_1218_),
    .S(_2621_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6601_ (.I(_2626_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6602_ (.I(_2620_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6603_ (.I0(_2610_),
    .I1(_1336_),
    .S(_2627_),
    .Z(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6604_ (.I(_2628_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6605_ (.I0(_2613_),
    .I1(_1633_),
    .S(_2627_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6606_ (.I(_2629_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6607_ (.I0(_2616_),
    .I1(_2081_),
    .S(_2627_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6608_ (.I(_2631_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6609_ (.I0(_2618_),
    .I1(_1548_),
    .S(_2627_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6610_ (.I(_2632_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6611_ (.A1(_2597_),
    .A2(_2559_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6612_ (.A1(_2561_),
    .A2(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6613_ (.I(_2634_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6614_ (.I0(_2596_),
    .I1(_0128_),
    .S(_2635_),
    .Z(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6615_ (.I(_2636_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6616_ (.I0(_2603_),
    .I1(_0256_),
    .S(_2635_),
    .Z(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6617_ (.I(_2638_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6618_ (.I0(_2605_),
    .I1(_0323_),
    .S(_2635_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6619_ (.I(_2639_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6620_ (.I0(_2608_),
    .I1(_0363_),
    .S(_2635_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6621_ (.I(_2640_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6622_ (.I(_2634_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6623_ (.I0(_2610_),
    .I1(_1695_),
    .S(_2641_),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6624_ (.I(_2642_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6625_ (.I0(_2613_),
    .I1(_1947_),
    .S(_2641_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6626_ (.I(_2643_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6627_ (.I0(_2616_),
    .I1(_2153_),
    .S(_2641_),
    .Z(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6628_ (.I(_2645_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6629_ (.I0(_2618_),
    .I1(_2152_),
    .S(_2641_),
    .Z(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6630_ (.I(_2646_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6631_ (.A1(_2582_),
    .A2(_2633_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6632_ (.I(_2647_),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6633_ (.I0(_2596_),
    .I1(_3209_),
    .S(_2648_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6634_ (.I(_2649_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6635_ (.I0(_2603_),
    .I1(_0252_),
    .S(_2648_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6636_ (.I(_2650_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6637_ (.I0(_2605_),
    .I1(_0403_),
    .S(_2648_),
    .Z(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6638_ (.I(_2652_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6639_ (.I0(_2608_),
    .I1(_0398_),
    .S(_2648_),
    .Z(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6640_ (.I(_2653_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6641_ (.I(_2647_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6642_ (.I0(_2610_),
    .I1(_1730_),
    .S(_2654_),
    .Z(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6643_ (.I(_2655_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6644_ (.I0(_2613_),
    .I1(_1971_),
    .S(_2654_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6645_ (.I(_2656_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6646_ (.I0(_2616_),
    .I1(_2173_),
    .S(_2654_),
    .Z(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6647_ (.I(_2658_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6648_ (.I0(_2618_),
    .I1(_2172_),
    .S(_2654_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6649_ (.I(_2659_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6650_ (.A1(net6),
    .A2(net5),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6651_ (.A1(_2561_),
    .A2(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6652_ (.I(_2661_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6653_ (.I0(_2558_),
    .I1(_1126_),
    .S(_2662_),
    .Z(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6654_ (.I(_2663_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6655_ (.I0(_2565_),
    .I1(_1122_),
    .S(_2662_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6656_ (.I(_2664_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6657_ (.I0(_2567_),
    .I1(_1463_),
    .S(_2662_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6658_ (.I(_2666_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6659_ (.I0(_2570_),
    .I1(_1579_),
    .S(_2662_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6660_ (.I(_2667_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6661_ (.I(_2661_),
    .Z(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6662_ (.I0(_2572_),
    .I1(_1593_),
    .S(_2668_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6663_ (.I(_2669_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6664_ (.I0(_2575_),
    .I1(_2055_),
    .S(_2668_),
    .Z(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6665_ (.I(_2670_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6666_ (.I0(_2578_),
    .I1(_1665_),
    .S(_2668_),
    .Z(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6667_ (.I(_2672_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6668_ (.I0(_2580_),
    .I1(_2313_),
    .S(_2668_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6669_ (.I(_2673_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6670_ (.A1(_2582_),
    .A2(_2660_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6671_ (.I(_2674_),
    .Z(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6672_ (.I0(_1295_),
    .I1(_2558_),
    .S(_2675_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6673_ (.I(_2676_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6674_ (.I0(_2710_),
    .I1(_2565_),
    .S(_2675_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6675_ (.I(_2677_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6676_ (.I0(_3092_),
    .I1(_2567_),
    .S(_2675_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6677_ (.I(_2679_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6678_ (.I0(_1546_),
    .I1(_2570_),
    .S(_2675_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6679_ (.I(_2680_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6680_ (.I(_2674_),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6681_ (.I0(_1627_),
    .I1(_2572_),
    .S(_2681_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6682_ (.I(_2682_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6683_ (.I0(_1917_),
    .I1(_2575_),
    .S(_2681_),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6684_ (.I(_2683_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6685_ (.I0(_1635_),
    .I1(_2578_),
    .S(_2681_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6686_ (.I(_2684_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6687_ (.I0(_2323_),
    .I1(_2580_),
    .S(_2681_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6688_ (.I(_2686_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6689_ (.D(_0000_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6690_ (.D(_0001_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6691_ (.D(_0002_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6692_ (.D(_0003_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6693_ (.D(_0004_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6694_ (.D(_0005_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6695_ (.D(_0006_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6696_ (.D(_0007_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6697_ (.D(_0008_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6698_ (.D(_0009_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6699_ (.D(_0010_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6700_ (.D(_0011_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6701_ (.D(_0012_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6702_ (.D(_0013_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6703_ (.D(_0014_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6704_ (.D(_0015_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6705_ (.D(_0016_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6706_ (.D(_0017_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6707_ (.D(_0018_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6708_ (.D(_0019_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6709_ (.D(_0020_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6710_ (.D(_0021_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6711_ (.D(_0022_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6712_ (.D(_0023_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6713_ (.D(_0024_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6714_ (.D(_0025_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6715_ (.D(_0026_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6716_ (.D(_0027_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6717_ (.D(_0028_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6718_ (.D(_0029_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6719_ (.D(_0030_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6720_ (.D(_0031_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.B[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6721_ (.D(_0032_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6722_ (.D(_0033_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6723_ (.D(_0034_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6724_ (.D(_0035_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6725_ (.D(_0036_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6726_ (.D(_0037_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6727_ (.D(_0038_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6728_ (.D(_0039_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6729_ (.D(_0040_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6730_ (.D(_0041_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6731_ (.D(_0042_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6732_ (.D(_0043_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6733_ (.D(_0044_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6734_ (.D(_0045_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6735_ (.D(_0046_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6736_ (.D(_0047_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6737_ (.D(_0048_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6738_ (.D(_0049_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6739_ (.D(_0050_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6740_ (.D(_0051_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6741_ (.D(_0052_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6742_ (.D(_0053_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6743_ (.D(_0054_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6744_ (.D(_0055_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6745_ (.D(_0056_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6746_ (.D(_0057_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6747_ (.D(_0058_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6748_ (.D(_0059_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6749_ (.D(_0060_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6750_ (.D(_0061_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6751_ (.D(_0062_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6752_ (.D(_0063_),
    .RN(net2),
    .CLK(net3),
    .Q(\k.A[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_178 (.Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_179 (.Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_180 (.Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_181 (.Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_182 (.Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_183 (.Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_184 (.Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_185 (.Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_186 (.Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_187 (.Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_188 (.Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_189 (.Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_190 (.Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_191 (.Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_192 (.Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__D (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_177 (.Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[22]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input2 (.I(io_in[23]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 input3 (.I(io_in[24]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[25]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[26]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[27]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[28]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[29]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(io_in[30]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(io_in[31]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(io_in[32]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(io_in[33]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(io_in[34]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(io_in[35]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(io_in[36]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(io_in[37]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output17 (.I(net17),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output18 (.I(net18),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output19 (.I(net19),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output20 (.I(net20),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output21 (.I(net21),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output22 (.I(net22),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output23 (.I(net23),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output24 (.I(net24),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output25 (.I(net25),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output26 (.I(net26),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output27 (.I(net27),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output28 (.I(net28),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output29 (.I(net29),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output30 (.I(net30),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output31 (.I(net31),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output32 (.I(net32),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output33 (.I(net33),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__D (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__D (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__D (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A2 (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A2 (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__I (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__I (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A1 (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A1 (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__B2 (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__B1 (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__B2 (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A2 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A2 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A1 (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__I (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__I (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__B2 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A1 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A2 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__A1 (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__B2 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__I (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__B2 (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A2 (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__B2 (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A1 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__A2 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A1 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__I (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A1 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A3 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A2 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__I (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A1 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__I (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__I1 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__B1 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A4 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__I (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__I (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__I (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A1 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A2 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__I (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A1 (.I(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A2 (.I(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A1 (.I(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__I (.I(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__I (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__B2 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A2 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__I (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A2 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__I (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A2 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__B2 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A2 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A3 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A1 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A2 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__I0 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A2 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__B1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__I (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__B1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A2 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A2 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A2 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A3 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A2 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A2 (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A1 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A2 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__I1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A4 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A3 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__I1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A4 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A3 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__I (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A3 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__B (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__I1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__I (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__I1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__I (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__I (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__I1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A3 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__I (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__I1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A2 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__B (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A3 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__B (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__B2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__B (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__B (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__I (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__B1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A3 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__I (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__I (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__I (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__I (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__I (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__B1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__I (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__I (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__I (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__I (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A4 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__B1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__I (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A3 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__B2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__I (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__I (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__I (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__B1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__B2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A3 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__B1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__B1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A3 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__I (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__B1 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__I (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__B2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A3 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A3 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__I (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__I (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A3 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A3 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A3 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__I (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__B1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__B1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__B1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__B1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__B2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__B1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__B1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__B1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A3 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__B2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__A1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__B2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__I (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__I (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__I (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__I (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__I (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A3 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A4 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__B1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__I (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__I1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__I (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A3 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__I (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A3 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__B (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__I (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A3 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__I0 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A4 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__I1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A4 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__B1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A3 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__B (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A3 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__B2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__B1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__I (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A3 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__I (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__I (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A3 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__I1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__I (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__I (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A1 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__B2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A3 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__I0 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__B2 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A2 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A3 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__I (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3364__I (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__I (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A2 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__I (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A3 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__B2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__B2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__C (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__I (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__C (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__C (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__B (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__I (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__I0 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A3 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__B2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__I (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__B2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__B2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__I (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A2 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3376__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__I (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A4 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__B1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__B1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A3 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A2 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__I1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A3 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__I (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__I (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__I1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__I (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__I (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__I0 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__I (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A2 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A2 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A2 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A2 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__I1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A3 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A3 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__B1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__B2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__B1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__I (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__B2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A2 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__B2 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__B1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__B2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A3 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__B1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A3 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__B1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__I0 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__B2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A4 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__B1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__B1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__I1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A3 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__B1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__B2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__B1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A3 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A4 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__B1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A3 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__I (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__I0 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__B2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__I1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__B1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A3 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A3 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A3 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__I (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__A1 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__I1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__B2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__B1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A1 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__I (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__B1 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__I (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__I (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__I (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__I (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__B2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__B2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__B1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__B2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__I (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__I0 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__I1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A3 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__I (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__B2 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A3 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__I1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__I (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__I0 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__I1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__I (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A3 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__C (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__I (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__C (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__C (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__C (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__C (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__B (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__I (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A4 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__B1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__A2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I0 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__I1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__I (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__I0 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A2 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__I1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__I0 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A3 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A3 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A2 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__B (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__B (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__I0 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__I1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__I0 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__I1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__I (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__I1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__I (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A3 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A3 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A3 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A3 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__B (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__B (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__I (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A3 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A3 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__B (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__B (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__B2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__I0 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A1 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__A2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__B (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A3 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__I0 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A2 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__I1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A1 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A1 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__I (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__I (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__I1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__I1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__I1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A2 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__I1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__I1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A3 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A3 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__I1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__I1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__B1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A1 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__I1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__I1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__B2 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__B2 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__B2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__B2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__A1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__C (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__C (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__C (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A2 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__B (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__B (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__I1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A2 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A2 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A2 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__I0 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A1 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A3 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__A2 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__I (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A2 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__I1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__I0 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A3 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__B1 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__B2 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__I (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A2 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__A2 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A2 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A1 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A2 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__B2 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A2 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__B (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__B (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__B (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__A2 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A2 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__C (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__B (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__B (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__B (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__I (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__B2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__B (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__I (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A3 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__B (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__B1 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__B2 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A1 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__I (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__I (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__I (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__B (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__B (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__I (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__B (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A3 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__I (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__B1 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A2 (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A3 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A2 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__I (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A2 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__I (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A3 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A3 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__B (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A3 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A3 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__B (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__I1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__I0 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__I1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__I1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__I (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__I (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__I1 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__I0 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__I1 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__I1 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__I1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__I0 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__I1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__I1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__I1 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__I0 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__I1 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__I1 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I1 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__I0 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__I1 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__I1 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__I1 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__I0 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__I1 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__I1 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__I (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__I1 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__I0 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__I1 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__I1 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__I1 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__I0 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__I1 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__I1 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__I (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__I (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__I (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__I0 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__I0 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__I0 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__I0 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__I (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__I (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__I0 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__I0 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__I0 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__I0 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__I0 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__I0 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__I0 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__I0 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__I0 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__I0 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__I0 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__I0 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__I0 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__I0 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__I0 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__I0 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__I0 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__I0 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__I0 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__I0 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__I0 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__I0 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__I0 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__I0 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__I0 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__I0 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__I0 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__I0 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__I (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__I (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__S (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__S (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__S (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__S (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__S (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__S (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__S (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__S (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__I (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__I (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__I (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__I (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__I (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__I (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__I (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__I (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__S (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__S (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__S (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__S (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__I (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__I (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__I (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__I (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__I (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__I (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__S (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__S (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__S (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__S (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A2 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__I (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A2 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A2 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A2 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A2 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__I (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__B1 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A2 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A2 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A1 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A1 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__I0 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A2 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__B2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__I (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A1 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A1 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A2 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A3 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A4 (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__B1 (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__I (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__I (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A4 (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__B1 (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A3 (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__I (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A2 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A2 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__I (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__I (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__B1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A2 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A2 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__I (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__B1 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__I (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__I (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A3 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__I (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__I (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__I (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A2 (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__I (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__I (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A4 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A2 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A2 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A2 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__I (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A2 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A1 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__I (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A1 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A2 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__I (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__I (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A2 (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__B1 (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__I (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__I (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A1 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__I (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A2 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A1 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A2 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A3 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A2 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__I (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__I (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A2 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A2 (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A2 (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A3 (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__B2 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A2 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__B2 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__I (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__B1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A3 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__I (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A1 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A1 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__I (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A1 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A1 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__I (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__B2 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__I (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A2 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A2 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__I (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A1 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__B1 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A2 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__I (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__I (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A3 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__I (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A4 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A2 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__I (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__I (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A2 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__I (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__I0 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A2 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A2 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B2 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A4 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__B1 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B1 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__I (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A2 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A1 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A1 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A3 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A2 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__B2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__B2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__B2 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A2 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A2 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A4 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__I (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A1 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A1 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A3 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A3 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__B2 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A1 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__I (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__I (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__I (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A1 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A1 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__I (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A1 (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A1 (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__B1 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A1 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__I (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__B2 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A1 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__B2 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A2 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__A1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__A1 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A1 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A1 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__A2 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__I (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__I (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__B1 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A2 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__I (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__B2 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A1 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A3 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A3 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A1 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A1 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A1 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__I (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A1 (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A1 (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__I (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A2 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A1 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A1 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A1 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A3 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A1 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A2 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A2 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A3 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A2 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A3 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A1 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A2 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__I (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__A2 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A2 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__I (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__I (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A1 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A1 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A4 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A4 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__I (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__I0 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__B1 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A2 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A2 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A2 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A3 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A2 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A3 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A1 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A2 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A2 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__I (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__I (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__B2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__I0 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__I (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A1 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A1 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__I1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A4 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__I1 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A2 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A2 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A1 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A1 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A1 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__B (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__I (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__B1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__B2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A2 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__B (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A1 (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__B (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__I (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__I (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__I0 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A1 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__I (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__I (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__I (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__B2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A2 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__I (.I(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A3 (.I(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__B (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A3 (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A1 (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A2 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__B (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__B (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A2 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__C (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A3 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__I (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__I1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__I (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__I (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__I (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__I (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A3 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__I (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__I (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A1 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__I (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__I (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__I (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__B2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__B2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__I (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__I (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__I (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A2 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A1 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__B2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A1 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__B2 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__B2 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__B2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__B2 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__I (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__B2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A3 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A2 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A2 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__I (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__I1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A2 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A3 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A2 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A1 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A2 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__I (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A2 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A2 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A2 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__I (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__I (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__I (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A2 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A1 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__I (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A1 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__I (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A2 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A1 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A1 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__I (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__B2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A1 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__I1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A2 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A2 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__I1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A2 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__B2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__I (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__B2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A2 (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A2 (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A2 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A2 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__B1 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__I (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__B1 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A1 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A1 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A3 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A1 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A2 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A1 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A1 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A2 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__I (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__I0 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__I (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A1 (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__I (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__I (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A2 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__I (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A2 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__I (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__B2 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__A1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__I (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__I (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A1 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__I (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A1 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__I (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__I (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__I (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__I (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A1 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A1 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A1 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A2 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__I (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__I (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__I (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__I (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__B1 (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A2 (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A2 (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__I (.I(\k.A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__I (.I(\k.A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A2 (.I(\k.A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__I (.I(\k.A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__I (.I(\k.A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A2 (.I(\k.A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A2 (.I(\k.A[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A2 (.I(\k.A[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A2 (.I(\k.A[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__I (.I(\k.A[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A2 (.I(\k.A[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A2 (.I(\k.A[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A1 (.I(\k.A[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__I (.I(\k.A[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A1 (.I(\k.A[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__I (.I(\k.A[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__I (.I(\k.A[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A1 (.I(\k.A[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A1 (.I(\k.A[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A2 (.I(\k.A[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A3 (.I(\k.A[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__I (.I(\k.A[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__I (.I(\k.A[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(\k.A[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A2 (.I(\k.A[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A4 (.I(\k.A[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__I (.I(\k.A[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(\k.A[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A1 (.I(\k.A[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__I (.I(\k.A[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__I (.I(\k.A[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__A2 (.I(\k.A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A1 (.I(\k.A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A1 (.I(\k.A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__I (.I(\k.A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A2 (.I(\k.A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__B2 (.I(\k.A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A1 (.I(\k.A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__I (.I(\k.A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A2 (.I(\k.A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__I (.I(\k.A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__I (.I(\k.A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A2 (.I(\k.A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A2 (.I(\k.A[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__I (.I(\k.A[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A2 (.I(\k.A[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__I (.I(\k.A[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(\k.A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(\k.A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__I (.I(\k.A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__I (.I(\k.A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(\k.A[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(\k.A[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__I (.I(\k.A[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__I (.I(\k.A[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I (.I(\k.A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__I (.I(\k.A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(\k.A[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__I (.I(\k.A[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A1 (.I(\k.A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__I (.I(\k.A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(\k.A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__I (.I(\k.A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(\k.A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A1 (.I(\k.A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__I (.I(\k.A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(\k.A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(\k.A[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__I (.I(\k.A[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__I (.I(\k.A[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(\k.A[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(\k.A[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__I (.I(\k.A[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(\k.A[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__I (.I(\k.A[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(\k.A[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__I (.I(\k.A[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I (.I(\k.A[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__I (.I(\k.A[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__I (.I(\k.A[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(\k.A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(\k.A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__I (.I(\k.A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A1 (.I(\k.A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__I (.I(\k.A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(\k.A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__I (.I(\k.B[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__I (.I(\k.B[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__I (.I(\k.B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__I (.I(\k.B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(\k.B[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__I (.I(\k.B[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(\k.B[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(\k.B[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(\k.B[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__I (.I(\k.B[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(\k.B[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__A2 (.I(\k.B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A2 (.I(\k.B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__I (.I(\k.B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3356__I (.I(\k.B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A1 (.I(\k.B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__I (.I(\k.B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A1 (.I(\k.B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__I (.I(\k.B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A1 (.I(\k.B[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__I (.I(\k.B[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A1 (.I(\k.B[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__I (.I(\k.B[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__I (.I(\k.B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__I (.I(\k.B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A1 (.I(\k.B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__I (.I(\k.B[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__I (.I(\k.B[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A2 (.I(\k.B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__I (.I(\k.B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__I (.I(\k.B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A2 (.I(\k.B[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__I (.I(\k.B[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__I (.I(\k.B[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A2 (.I(\k.B[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(\k.B[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__I (.I(\k.B[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(\k.B[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(\k.B[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__I (.I(\k.B[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__I (.I(\k.B[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A2 (.I(\k.B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A2 (.I(\k.B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__I (.I(\k.B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__I (.I(\k.B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net34;
 assign io_oeb[10] = net44;
 assign io_oeb[11] = net45;
 assign io_oeb[12] = net46;
 assign io_oeb[13] = net47;
 assign io_oeb[14] = net48;
 assign io_oeb[15] = net49;
 assign io_oeb[16] = net50;
 assign io_oeb[17] = net51;
 assign io_oeb[18] = net52;
 assign io_oeb[19] = net53;
 assign io_oeb[1] = net35;
 assign io_oeb[20] = net54;
 assign io_oeb[21] = net55;
 assign io_oeb[22] = net177;
 assign io_oeb[23] = net178;
 assign io_oeb[24] = net179;
 assign io_oeb[25] = net180;
 assign io_oeb[26] = net181;
 assign io_oeb[27] = net182;
 assign io_oeb[28] = net183;
 assign io_oeb[29] = net184;
 assign io_oeb[2] = net36;
 assign io_oeb[30] = net185;
 assign io_oeb[31] = net186;
 assign io_oeb[32] = net187;
 assign io_oeb[33] = net188;
 assign io_oeb[34] = net189;
 assign io_oeb[35] = net190;
 assign io_oeb[36] = net191;
 assign io_oeb[37] = net192;
 assign io_oeb[3] = net37;
 assign io_oeb[4] = net38;
 assign io_oeb[5] = net39;
 assign io_oeb[6] = net40;
 assign io_oeb[7] = net41;
 assign io_oeb[8] = net42;
 assign io_oeb[9] = net43;
 assign io_out[0] = net56;
 assign io_out[1] = net57;
 assign io_out[22] = net61;
 assign io_out[23] = net62;
 assign io_out[24] = net63;
 assign io_out[25] = net64;
 assign io_out[26] = net65;
 assign io_out[27] = net66;
 assign io_out[28] = net67;
 assign io_out[29] = net68;
 assign io_out[2] = net58;
 assign io_out[30] = net69;
 assign io_out[31] = net70;
 assign io_out[32] = net71;
 assign io_out[33] = net72;
 assign io_out[34] = net73;
 assign io_out[35] = net74;
 assign io_out[36] = net75;
 assign io_out[37] = net76;
 assign io_out[3] = net59;
 assign io_out[4] = net60;
 assign la_data_out[0] = net77;
 assign la_data_out[10] = net87;
 assign la_data_out[11] = net88;
 assign la_data_out[12] = net89;
 assign la_data_out[13] = net90;
 assign la_data_out[14] = net91;
 assign la_data_out[15] = net92;
 assign la_data_out[16] = net93;
 assign la_data_out[17] = net94;
 assign la_data_out[18] = net95;
 assign la_data_out[19] = net96;
 assign la_data_out[1] = net78;
 assign la_data_out[20] = net97;
 assign la_data_out[21] = net98;
 assign la_data_out[22] = net99;
 assign la_data_out[23] = net100;
 assign la_data_out[24] = net101;
 assign la_data_out[25] = net102;
 assign la_data_out[26] = net103;
 assign la_data_out[27] = net104;
 assign la_data_out[28] = net105;
 assign la_data_out[29] = net106;
 assign la_data_out[2] = net79;
 assign la_data_out[30] = net107;
 assign la_data_out[31] = net108;
 assign la_data_out[32] = net109;
 assign la_data_out[33] = net110;
 assign la_data_out[34] = net111;
 assign la_data_out[35] = net112;
 assign la_data_out[36] = net113;
 assign la_data_out[37] = net114;
 assign la_data_out[38] = net115;
 assign la_data_out[39] = net116;
 assign la_data_out[3] = net80;
 assign la_data_out[40] = net117;
 assign la_data_out[41] = net118;
 assign la_data_out[42] = net119;
 assign la_data_out[43] = net120;
 assign la_data_out[44] = net121;
 assign la_data_out[45] = net122;
 assign la_data_out[46] = net123;
 assign la_data_out[47] = net124;
 assign la_data_out[48] = net125;
 assign la_data_out[49] = net126;
 assign la_data_out[4] = net81;
 assign la_data_out[50] = net127;
 assign la_data_out[51] = net128;
 assign la_data_out[52] = net129;
 assign la_data_out[53] = net130;
 assign la_data_out[54] = net131;
 assign la_data_out[55] = net132;
 assign la_data_out[56] = net133;
 assign la_data_out[57] = net134;
 assign la_data_out[58] = net135;
 assign la_data_out[59] = net136;
 assign la_data_out[5] = net82;
 assign la_data_out[60] = net137;
 assign la_data_out[61] = net138;
 assign la_data_out[62] = net139;
 assign la_data_out[63] = net140;
 assign la_data_out[6] = net83;
 assign la_data_out[7] = net84;
 assign la_data_out[8] = net85;
 assign la_data_out[9] = net86;
 assign user_irq[0] = net141;
 assign user_irq[1] = net142;
 assign user_irq[2] = net143;
 assign wbs_ack_o = net144;
 assign wbs_dat_o[0] = net145;
 assign wbs_dat_o[10] = net155;
 assign wbs_dat_o[11] = net156;
 assign wbs_dat_o[12] = net157;
 assign wbs_dat_o[13] = net158;
 assign wbs_dat_o[14] = net159;
 assign wbs_dat_o[15] = net160;
 assign wbs_dat_o[16] = net161;
 assign wbs_dat_o[17] = net162;
 assign wbs_dat_o[18] = net163;
 assign wbs_dat_o[19] = net164;
 assign wbs_dat_o[1] = net146;
 assign wbs_dat_o[20] = net165;
 assign wbs_dat_o[21] = net166;
 assign wbs_dat_o[22] = net167;
 assign wbs_dat_o[23] = net168;
 assign wbs_dat_o[24] = net169;
 assign wbs_dat_o[25] = net170;
 assign wbs_dat_o[26] = net171;
 assign wbs_dat_o[27] = net172;
 assign wbs_dat_o[28] = net173;
 assign wbs_dat_o[29] = net174;
 assign wbs_dat_o[2] = net147;
 assign wbs_dat_o[30] = net175;
 assign wbs_dat_o[31] = net176;
 assign wbs_dat_o[3] = net148;
 assign wbs_dat_o[4] = net149;
 assign wbs_dat_o[5] = net150;
 assign wbs_dat_o[6] = net151;
 assign wbs_dat_o[7] = net152;
 assign wbs_dat_o[8] = net153;
 assign wbs_dat_o[9] = net154;
endmodule

