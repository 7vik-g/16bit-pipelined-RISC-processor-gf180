* NGSPICE file created from processor.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

.subckt processor Dataw_en Serial_input Serial_output clk data_mem_addr[0] data_mem_addr[1]
+ data_mem_addr[2] data_mem_addr[3] data_mem_addr[4] data_mem_addr[5] data_mem_addr[6]
+ data_mem_addr[7] hlt instr[0] instr[10] instr[11] instr[12] instr[13] instr[14]
+ instr[15] instr[1] instr[2] instr[3] instr[4] instr[5] instr[6] instr[7] instr[8]
+ instr[9] instr_mem_addr[0] instr_mem_addr[10] instr_mem_addr[11] instr_mem_addr[12]
+ instr_mem_addr[1] instr_mem_addr[2] instr_mem_addr[3] instr_mem_addr[4] instr_mem_addr[5]
+ instr_mem_addr[6] instr_mem_addr[7] instr_mem_addr[8] instr_mem_addr[9] read_data[0]
+ read_data[10] read_data[11] read_data[12] read_data[13] read_data[14] read_data[15]
+ read_data[1] read_data[2] read_data[3] read_data[4] read_data[5] read_data[6] read_data[7]
+ read_data[8] read_data[9] reset start vdd vss write_data[0] write_data[10] write_data[11]
+ write_data[12] write_data[13] write_data[14] write_data[15] write_data[1] write_data[2]
+ write_data[3] write_data[4] write_data[5] write_data[6] write_data[7] write_data[8]
+ write_data[9]
XFILLER_228_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3140__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3155_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3086_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_227_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5160__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2953__I _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__RN net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_243_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3988_ _0882_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4878__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2939_ net49 _0765_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_206_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2954__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4609_ _1923_ _1954_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5188__RN net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2890__B1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2863__I Arithmetic_Logic_Unit.ALU_001.p_Z vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4631__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5112__RN net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3694__I _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2945__A1 Control_unit1.instr_stage1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5179__RN net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5033__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3122__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5183__CLK clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout260_I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _0122_ net344 clknet_leaf_46_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_188_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4622__A1 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3911_ _1160_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4891_ net3 net123 clknet_leaf_9_clk Control_unit1.instr_stage1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3842_ _1303_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3189__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3773_ _1352_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2724_ _0573_ _0579_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2655_ _2337_ _2137_ _2138_ _2318_ _2339_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ _0536_ net321 clknet_leaf_51_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2586_ _2249_ _2263_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4917__RN net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2948__I _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4325_ _1659_ _1753_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout105 net107 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout116 net117 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout127 net128 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout138 net140 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout149 net150 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ _1603_ _1705_ _1709_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3113__A1 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3207_ _0970_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4187_ _1627_ _1664_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3138_ _2363_ _0584_ _0911_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_216_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3069_ _0865_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3416__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5056__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3019__I _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3352__A1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3104__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__RN net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2593__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3591__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2440_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout106_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3343__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3894__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4110_ _1585_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5090_ _0252_ net101 clknet_leaf_110_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4041_ _1503_ _1560_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_204_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3646__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4943_ _0105_ net342 clknet_leaf_46_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_212_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4071__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5079__CLK clknet_leaf_102_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4874_ Control_unit1.instr_stage1\[9\] net129 clknet_leaf_4_clk Control_unit2.instr_stage2\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3825_ _1348_ _1408_ _1413_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3756_ _1312_ _1367_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3582__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2707_ _2161_ _2365_ _0566_ _2164_ _2208_ _2337_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3687_ _1150_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2638_ _2317_ _2096_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4916__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5357_ _0519_ net311 clknet_leaf_50_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2569_ _2108_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3885__A2 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _1745_ _1739_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5288_ _0450_ net187 clknet_leaf_66_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_210_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4239_ _1696_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_227_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3573__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3972__I _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3325__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2588__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__A2 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5221__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5371__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3610_ _1191_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout223_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4939__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _1900_ _1937_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ net19 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3472_ _1159_ _1154_ _1162_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _0373_ net175 clknet_leaf_92_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2423_ net37 net1 _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3867__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5142_ _0304_ net158 clknet_leaf_95_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5073_ _0235_ net180 clknet_leaf_104_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_211_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_84_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4024_ _1482_ _1551_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_225_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_99_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4044__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2961__I _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4926_ _0088_ net341 clknet_leaf_45_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ Stack_pointer.SP_next\[1\] net115 clknet_leaf_8_clk Stack_pointer.SP\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_205_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clk_I clknet_4_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _1321_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4788_ _2067_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3555__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3739_ _1195_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_37_clk_I clknet_4_13_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3307__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2530__A2 Arithmetic_Logic_Unit.ALU_001.Y_CY\[4\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4128__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3967__I _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3546__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3207__I _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4274__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout173_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout340_I net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2972_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_188_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4711_ _2005_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _1910_ _1971_ _1975_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3537__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5117__CLK clknet_leaf_90_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4573_ _1929_ _1930_ _1932_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4501__I _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3524_ _0794_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_200_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3455_ _1145_ _1136_ _1148_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2406_ Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\] _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3386_ _0962_ _1098_ _1101_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2956__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5125_ _0287_ net174 clknet_leaf_100_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5056_ _0218_ net244 clknet_leaf_78_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4265__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4007_ _1459_ _1538_ _1541_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_226_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3787__I _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4909_ _0071_ net346 clknet_leaf_43_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_205_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3528__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4411__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2751__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output67_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4256__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4008__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3519__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4321__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3240_ _0996_ _0984_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2776__I _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout290_I net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3171_ _0802_ _0944_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3058__I0 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2955_ _2144_ _0779_ _0784_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2886_ net79 _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _1951_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4556_ _1916_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3507_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4487_ _1866_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3438_ _1045_ _1128_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2686__I _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3369_ _1060_ _1084_ _1089_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _0270_ net162 clknet_leaf_98_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5039_ _0201_ net254 clknet_leaf_76_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3997__A1 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3049__I0 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4410__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2421__A1 Control_unit1.instr_stage1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_114_clk clknet_4_0_0_clk clknet_leaf_114_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput42 net42 data_mem_addr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_218_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput53 net53 instr_mem_addr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput64 net64 write_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput75 net75 write_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_235_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4477__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2488__A1 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4229__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4316__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2660__A1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2740_ _0577_ _0582_ _0583_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA_fanout136_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_105_clk clknet_4_9_0_clk clknet_leaf_105_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2671_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3 _2108_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout303_I net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__A1 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _1735_ _1812_ _1818_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5390_ _0552_ net322 clknet_leaf_52_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4341_ net23 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout309 net313 net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4272_ _1621_ _1717_ _1719_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3223_ _0797_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3140__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3154_ _0931_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5305__CLK clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3085_ _0700_ _0701_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_236_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4640__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4226__I _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3987_ _1491_ _1522_ _1527_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_241_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2938_ net50 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_206_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2869_ net70 _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4608_ _1864_ _1952_ _1955_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4539_ _1902_ _1903_ _1906_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3305__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2890__A1 Control_unit2.instr_stage2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2890__B2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4136__I _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4871__RN net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3975__I _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4822__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4972__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3215__I _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3122__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4046__I _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3910_ _1324_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout253_I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4890_ net17 net116 clknet_leaf_8_clk Control_unit1.instr_stage1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__A1 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3841_ _1418_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4386__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3772_ _1379_ _1372_ _1380_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_207_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2723_ _0561_ _0562_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ _2082_ _2338_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5373_ _0535_ net321 clknet_leaf_50_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2585_ _2272_ _2207_ _2252_ _2273_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4324_ _1328_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout106 net108 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout117 net118 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_236_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout128 net129 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout139 net140 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ _1604_ _1706_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3206_ _0967_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4186_ _1621_ _1663_ _1665_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_210_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2964__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3137_ _2203_ _2294_ _0914_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3068_ _2106_ _0601_ _2252_ _0612_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4853__RN net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__CLK clknet_leaf_119_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4301__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5097__RN net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5000__CLK clknet_leaf_63_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5150__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3343__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5021__RN net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4040_ _1449_ _1558_ _1562_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4868__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2784__I _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4942_ _0104_ net342 clknet_leaf_47_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2606__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4835__RN net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4873_ Control_unit1.instr_stage1\[8\] net129 clknet_leaf_4_clk Control_unit2.instr_stage2\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3824_ _1349_ _1409_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_242_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3031__A1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3755_ _1307_ _1366_ _1369_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2706_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_203_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3686_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2637_ _2281_ _2258_ _2308_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3056__S _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3334__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5356_ _0518_ net275 clknet_leaf_60_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2568_ _2141_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4307_ net30 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _0449_ net192 clknet_leaf_69_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2499_ _2184_ _2110_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4238_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3098__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I read_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4169_ _1607_ _1650_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_94_clk clknet_4_8_0_clk clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_210_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5023__CLK clknet_leaf_55_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__RN net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5173__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4770__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3325__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4522__A1 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2836__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_85_clk clknet_4_10_0_clk clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4324__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3540_ _1159_ _1211_ _1214_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout216_I net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__RN net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3471_ _1161_ _1157_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _0372_ net170 clknet_leaf_94_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2422_ _2114_ Control_unit1.instr_stage1\[2\] _2115_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4513__A1 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _0303_ net174 clknet_leaf_100_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_233_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5072_ _0234_ net246 clknet_leaf_79_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4023_ _1532_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2827__A1 Control_unit1.instr_stage1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3403__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5046__CLK clknet_leaf_102_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_76_clk clknet_4_14_0_clk clknet_leaf_76_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__RN net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4925_ _0087_ net340 clknet_leaf_47_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5196__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4856_ Stack_pointer.SP_next\[0\] net122 clknet_leaf_9_clk Stack_pointer.SP\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3807_ _1390_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4787_ _2058_ net51 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4752__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3555__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3738_ _1285_ _1353_ _1357_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3669_ _1300_ _1289_ _1301_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4504__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5339_ _0501_ net305 clknet_leaf_58_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_67_clk clknet_4_9_0_clk clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_244_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_244_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4144__I _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4743__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__RN net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2809__A1 Control_unit1.instr_stage1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3223__I _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_58_clk clknet_4_12_0_clk clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_187_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4906__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2971_ net28 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout333_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4710_ _0994_ _2013_ _2018_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4641_ _1911_ _1972_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3893__I _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4572_ _1878_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3523_ _1134_ _1189_ _1203_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3454_ _1147_ _1139_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ _2083_ _2097_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3385_ _1037_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _0286_ net86 clknet_leaf_116_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout79_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5055_ _0217_ net244 clknet_leaf_78_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_49_clk clknet_4_15_0_clk clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_211_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4006_ _1460_ _1539_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2972__I _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3225__A1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4908_ _0070_ net333 clknet_leaf_41_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3776__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4839_ _0041_ net148 clknet_leaf_18_clk net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4725__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5206__RN net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5211__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2503__A3 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5361__CLK clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4139__I _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4929__CLK clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3978__I _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2882__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3216__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4716__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_83_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4192__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3218__I _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_98_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3170_ _0795_ _0943_ _0945_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout283_I net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_21_clk_I clknet_4_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3455__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_36_clk_I clknet_4_13_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3058__I1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2954_ _0781_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2430__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2885_ net54 _0716_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4707__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _1887_ _1959_ _1964_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ net18 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3506_ net18 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4486_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5384__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3437_ _0979_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3064__S _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_109_clk_I clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3368_ _1011_ _1085_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _0269_ net90 clknet_leaf_114_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3299_ _0977_ _1036_ _1044_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _0200_ net254 clknet_leaf_75_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input11_I instr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3049__I1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2421__A2 Control_unit1.instr_stage1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__I _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4174__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput43 net43 data_mem_addr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput54 net54 instr_mem_addr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput65 net65 write_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5107__CLK clknet_leaf_114_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2660__A2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2670_ _2354_ net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout129_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4165__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3912__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ _1343_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4271_ _1623_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3222_ _0968_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input3_I instr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3153_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3140__A3 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3084_ _2119_ _2087_ _0880_ _2085_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4507__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ _1492_ _1523_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_241_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2937_ _0722_ _0764_ _0767_ _0750_ _0768_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_221_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2868_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4607_ _1919_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2799_ Control_unit1.instr_stage1\[6\] _0630_ _0631_ _0650_ _0651_ _0652_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4538_ _1904_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3903__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4469_ _1755_ _1852_ _1855_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_232_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3419__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4395__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_220_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_210_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3991__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4327__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2633__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout246_I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3840_ _1416_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4386__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _1331_ _1373_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2722_ _2375_ _0579_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_160_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4138__A2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2653_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_218_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2584_ _2230_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5372_ _0534_ net310 clknet_leaf_60_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _1755_ _1751_ _1757_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout118 net128 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout129 net153 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4254_ _1600_ _1705_ _1708_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3205_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4185_ _1623_ _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3136_ _2158_ _2183_ _2229_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_132_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4237__I _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3067_ _2234_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2624__A2 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2980__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3969_ _1468_ _1514_ _1516_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4129__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4301__A2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4147__I _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3051__I _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2615__A2 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3879__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout196_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4941_ _0103_ net340 clknet_leaf_47_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3896__I _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4872_ Control_unit1.instr_stage1\[7\] net124 clknet_leaf_10_clk Control_unit2.instr_stage2\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_221_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3823_ _1344_ _1408_ _1412_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_242_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3754_ _1308_ _1367_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2705_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[13\].i3 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3685_ _2296_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4520__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2636_ _2322_ net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _0517_ net309 clknet_leaf_60_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2567_ _2256_ net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2542__A1 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4306_ _1310_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5286_ _0448_ net185 clknet_leaf_106_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2498_ _2190_ net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4812__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4237_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3098__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4168_ _1603_ _1649_ _1653_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3119_ _0822_ _0899_ _0904_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4099_ _1601_ _1598_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4962__CLK clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4598__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2924__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5318__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_221_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__A2 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2781__A1 Stack_pointer.SP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2836__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_235_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4038__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3013__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__A1 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4340__I _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2772__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout111_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout209_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3470_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2421_ Control_unit1.instr_stage1\[3\] Control_unit1.instr_stage1\[1\] _2116_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4835__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5140_ _0302_ net86 clknet_leaf_116_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5071_ _0233_ net246 clknet_leaf_79_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_211_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4985__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4022_ _1530_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2827__A2 Control_unit1.instr_stage1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4515__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _0086_ net332 clknet_leaf_40_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4855_ _0057_ net349 clknet_leaf_44_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_221_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3806_ _1388_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4786_ _2058_ net76 net52 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3737_ _1354_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4250__I _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3668_ _1202_ _1291_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4992__RN net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2619_ _2131_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4504__A2 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3599_ _1176_ _1252_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5338_ _0500_ net273 clknet_leaf_62_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_27_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4268__A1 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ _0431_ net185 clknet_leaf_106_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3491__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5140__CLK clknet_leaf_116_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4160__I _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4983__RN net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2506__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3504__I _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout290 net302 net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2970_ _0778_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2993__A1 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout326_I net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4640_ _1907_ _1971_ _1974_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4571_ _1920_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3522_ _1202_ _1193_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3453_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5013__CLK clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2404_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3384_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3170__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ _0285_ net84 clknet_leaf_116_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_217_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3414__I _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5054_ _0216_ net244 clknet_leaf_78_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5163__CLK clknet_leaf_89_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4005_ _1507_ _1538_ _1540_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__A1 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _0069_ net335 clknet_leaf_42_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4838_ _0040_ net149 clknet_leaf_18_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[0\].i2
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_72_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4725__A2 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _1019_ _2052_ _2055_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3161__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4661__A1 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4413__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2975__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5036__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4956__RN net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5186__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3234__I _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4652__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__RN net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4065__I _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2953_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2966__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2884_ _0710_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ _1888_ _1960_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4554_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3391__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3505_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4485_ _1724_ _1286_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout91_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3436_ _1132_ _1126_ _1133_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3143__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3367_ _1009_ _1084_ _1088_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5372__RN net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _0268_ net90 clknet_leaf_114_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3298_ _1043_ _1039_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5037_ _0199_ net250 clknet_leaf_75_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5124__RN net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5059__CLK clknet_leaf_110_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput44 net44 data_mem_addr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput55 net79 instr_mem_addr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output72_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput66 net66 write_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3134__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5363__RN net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2893__I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5115__RN net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_201_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3229__I _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4270_ _1699_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3221_ _0980_ _0969_ _0981_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3152_ _2089_ _0701_ _0881_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_6590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3083_ _0687_ Control_unit2.instr_decoder2.A\[1\] _2140_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_236_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5201__CLK clknet_leaf_114_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3985_ _1488_ _1522_ _1526_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_225_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2939__A1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ net49 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3600__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2867_ _2088_ _0703_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5351__CLK clknet_leaf_64_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4606_ _1953_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4919__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2798_ Stack_pointer.SP\[3\] _0632_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4537_ _1868_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4468_ _1756_ _1853_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3116__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3419_ _1025_ _1118_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4399_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3419__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_82_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_97_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_35_clk_I clknet_4_13_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3512__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5224__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout141_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_108_clk_I clknet_4_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3770_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout239_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3594__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2721_ _0573_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_203_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2652_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_199_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3346__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _0533_ net309 clknet_leaf_60_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2583_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _1756_ _1753_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout119 net121 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4253_ _1601_ _1706_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_234_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3204_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ _1639_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3135_ _2129_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4518__I _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3066_ _0687_ _2234_ Control_unit2.instr_decoder2.A\[2\] Control_unit2.instr_decoder2.A\[1\]
+ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_243_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4074__A2 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3821__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3968_ _1470_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ _2088_ _0703_ _0705_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3899_ _1462_ _1455_ _1464_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4891__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5247__CLK clknet_leaf_77_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3507__I _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3879__A2 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5309__RN net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3500__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3242__I _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout189_I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ _0102_ net311 clknet_leaf_50_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3803__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ Control_unit1.instr_stage1\[6\] net124 clknet_leaf_10_clk Control_unit2.instr_stage2\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_209_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3822_ _1345_ _1409_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3567__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3753_ _1365_ _1366_ _1368_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2704_ _0560_ _0563_ _2278_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3684_ _1311_ _1302_ _1313_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2635_ _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5354_ _0516_ net275 clknet_leaf_60_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_173_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2566_ _2255_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4305_ _1741_ _1737_ _1743_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ _0447_ net185 clknet_leaf_106_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2497_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4236_ _0883_ _0964_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4167_ _1604_ _1650_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3118_ _0824_ _0900_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4098_ _1142_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2991__I _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3049_ _0812_ _2282_ _0851_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_227_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_221_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3558__A1 Control_unit2.instr_stage2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4711__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3327__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4038__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2406__I Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout90 net91 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2772__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3237__I _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2420_ net77 net78 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout104_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5070_ _0232_ net242 clknet_leaf_80_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_215_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4277__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ _1520_ _1544_ _1549_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_238_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4029__A2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3788__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4923_ _0085_ net329 clknet_leaf_39_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_209_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_221_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4854_ _0056_ net349 clknet_leaf_45_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_222_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3805_ _1315_ _1396_ _1401_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4785_ net52 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4201__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4531__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5092__CLK clknet_leaf_103_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3736_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2763__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3667_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2618_ _2152_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3598_ _1168_ _1251_ _1253_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5337_ _0499_ net305 clknet_leaf_60_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2549_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3 _2109_ _2238_ _2149_ _2239_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_216_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5268_ _0430_ net104 clknet_leaf_118_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input34_I reset vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4268__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ _1609_ _1684_ _1686_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _0361_ net226 clknet_leaf_84_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_217_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__A2 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3951__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2506__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout280 net303 net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout291 net295 net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4616__I _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3520__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4351__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout319_I net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4570_ _1917_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3521_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3452_ net30 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2403_ _2078_ _2081_ Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\] _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3383_ _1096_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ _0284_ net84 clknet_leaf_115_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5308__CLK clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5053_ _0215_ net243 clknet_leaf_81_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_242_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4004_ _1456_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_226_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ _0068_ net334 clknet_leaf_42_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2433__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4837_ _0039_ net149 clknet_leaf_33_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[14\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4768_ _0831_ _2053_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2736__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3719_ _1341_ _1337_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4699_ _1927_ _2008_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2672__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3340__I _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_117_clk clknet_4_1_0_clk clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4171__I _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4975__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3152__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout171_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3250__I _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout269_I net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4404__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2952_ _0777_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_108_clk clknet_4_1_0_clk clknet_leaf_108_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2883_ _0708_ _0711_ _0718_ _0720_ _0721_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ _1884_ _1959_ _1963_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_198_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4553_ _1916_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3504_ _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4484_ _2143_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3435_ _1043_ _1128_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5130__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3143__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3366_ _1058_ _1085_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _0267_ net162 clknet_leaf_98_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3297_ _0788_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5280__CLK clknet_leaf_76_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ _0198_ net239 clknet_leaf_73_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2485__B _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4848__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4643__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4998__CLK clknet_leaf_63_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4159__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput45 net45 data_mem_addr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput56 net56 instr_mem_addr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput67 net67 write_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output65_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4874__RN net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4398__A1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5003__CLK clknet_leaf_57_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_9_clk_I clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5153__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3373__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3245__I _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3125__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3220_ _0792_ _0971_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3151_ _0930_ Control_unit2.instr_stage2\[9\] Control_unit2.instr_stage2\[10\] _0931_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3082_ _0747_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_5890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4865__RN net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ _1489_ _1523_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_206_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2935_ _0701_ _0748_ _0714_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_241_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2866_ _2089_ _0704_ Arithmetic_Logic_Unit.ALU_001.p_Z _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _1950_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2797_ Stack_pointer.SP\[3\] _0642_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4561__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4536_ net21 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3155__I _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _1750_ _1852_ _1854_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3418_ _1020_ _1117_ _1120_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4398_ _1724_ _1226_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2994__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3349_ _0980_ _1071_ _1077_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _0181_ net306 clknet_leaf_57_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__CLK clknet_leaf_118_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4856__RN net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5176__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2563__B1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4791__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2720_ _0577_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_fanout134_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__RN net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2651_ _2336_ net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_172_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout301_I net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5024__RN net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2582_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[7\].i3 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5370_ _0532_ net309 clknet_leaf_60_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ net33 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4252_ _1648_ _1705_ _1707_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout109 net110 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3203_ _0964_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4183_ _1636_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3703__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5049__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3134_ _0687_ _0601_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3065_ _0863_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3282__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5199__CLK clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4534__I _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3967_ _1498_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4782__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2918_ Control_unit2.instr_stage2\[9\] _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_30_clk clknet_4_6_0_clk clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3898_ _1463_ _1457_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2989__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2849_ Control_unit2.instr_stage2\[4\] _0681_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3337__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4519_ _1866_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_97_clk clknet_4_8_0_clk clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__RN net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_187_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_21_clk clknet_4_3_0_clk clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3328__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5006__RN net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_88_clk clknet_4_10_0_clk clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3500__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5341__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4909__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout251_I net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_206_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4870_ Control_unit1.instr_stage1\[5\] net125 clknet_leaf_9_clk Control_unit2.instr_stage2\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout349_I net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3016__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3821_ _1340_ _1408_ _1411_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3752_ _1303_ _1367_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_clk clknet_4_4_0_clk clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_203_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2703_ _0561_ _0562_ _2375_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3683_ _1312_ _1304_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3319__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4516__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_81_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2634_ _2316_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2565_ _2234_ _2248_ _2254_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5353_ _0515_ net309 clknet_leaf_60_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_154_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4304_ _1742_ _1739_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2496_ _2188_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5284_ _0446_ net104 clknet_leaf_118_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_clkbuf_leaf_96_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4235_ _1632_ _1690_ _1695_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_79_clk clknet_4_11_0_clk clknet_leaf_79_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_190_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4166_ _1600_ _1649_ _1652_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3117_ _2354_ _0899_ _0903_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4097_ _1306_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3048_ _0854_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_34_clk_I clknet_4_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3007__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _0161_ net273 clknet_leaf_63_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_212_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3558__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2512__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[4\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_49_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3730__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5364__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_107_clk_I clknet_4_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4746__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5227__RN net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net82 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_243_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout91 net92 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_168_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_6_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2524__A3 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout299_I net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ _1478_ _1545_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_1_clk clknet_4_1_0_clk clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_238_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4881__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ _0084_ net333 clknet_leaf_41_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_212_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4853_ _0055_ net348 clknet_leaf_43_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2460__A2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4737__A1 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3804_ _1316_ _1397_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__CLK clknet_leaf_104_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4784_ _2063_ _0731_ _2066_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3735_ _1351_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3428__I _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3960__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3666_ _2211_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2617_ _2281_ _2235_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3597_ _1171_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5336_ _0498_ net263 clknet_leaf_64_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2548_ _2130_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4259__I _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5267_ _0429_ net96 clknet_leaf_117_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2479_ _2113_ _2155_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ _1611_ _1685_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5198_ _0360_ net223 clknet_leaf_83_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input27_I read_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4149_ _1638_ _1640_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3779__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4722__I _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A1 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3400__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3338__I _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3951__A2 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3467__A1 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout270 net280 net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout281 net283 net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout292 net294 net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_212_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4719__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3520_ net27 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout214_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3451_ _0990_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2402_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[0\].i3 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3382_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5121_ _0283_ net161 clknet_leaf_98_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4079__I _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5052_ _0214_ net234 clknet_leaf_71_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4003_ _1532_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3711__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4905_ _0067_ net334 clknet_leaf_42_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_240_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2433__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3630__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4836_ _0038_ net284 clknet_leaf_33_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[13\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4186__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3158__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _1013_ _2052_ _2054_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3933__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3718_ _1175_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4698_ _0976_ _2006_ _2011_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3649_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5319_ _0481_ net263 clknet_leaf_65_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3449__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2672__A2 Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3621__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_236_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_223_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3924__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_197_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3152__A3 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_212_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5082__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout164_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2951_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3612__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout331_I net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4362__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2882_ net54 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4621_ _1885_ _1960_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4168__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4552_ _1724_ _1033_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3915__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3503_ _1031_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3706__I _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4483_ _1773_ _1858_ _1863_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3434_ _0976_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3365_ _1005_ _1084_ _1087_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5104_ _0266_ net246 clknet_leaf_79_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_246_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3296_ _0974_ _1036_ _1042_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4537__I _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ _0197_ net306 clknet_leaf_57_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3441__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2654__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3603__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4819_ _0021_ net346 clknet_leaf_42_clk net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_clkbuf_4_14_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput46 net46 hlt vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput57 net57 instr_mem_addr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput68 net68 write_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output58_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3351__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4942__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4398__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3526__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_234_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3150_ Control_unit2.instr_stage2\[8\] _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_6570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout281_I net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3081_ Control_unit2.instr_stage2\[9\] Control_unit2.instr_stage2\[10\] _0878_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3261__I _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3983_ _1485_ _1522_ _1525_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4092__I _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2934_ net49 _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_206_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2865_ Control_unit2.instr_stage2\[11\] _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4604_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2796_ Stack_pointer.SP\[3\] _0621_ _0635_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4535_ _1866_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2572__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4466_ _1752_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3417_ _1021_ _1118_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4313__A2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _1773_ _1804_ _1809_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3348_ _1045_ _1073_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3279_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _0180_ net236 clknet_leaf_57_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2627__A2 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2515__I _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4001__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2563__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2563__B2 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4177__I _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3815__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5120__CLK clknet_leaf_86_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4791__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2650_ _2335_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout127_I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5270__CLK clknet_leaf_106_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2581_ _2268_ _2269_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2554__A1 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _1324_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4251_ _1597_ _1706_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3202_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4988__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4182_ _1661_ _1655_ _1662_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input1_I Serial_input vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3133_ _2242_ _2247_ _2268_ _2269_ _0912_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3064_ _0838_ _0612_ _0850_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_209_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3282__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3966_ _1495_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2917_ net59 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3897_ _1146_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2793__A1 Stack_pointer.SP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2848_ _0690_ _0691_ net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2779_ Stack_pointer.SP\[0\] _0621_ _0629_ _0634_ Stack_pointer.SP_next\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4518_ _2321_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4449_ _1731_ _1839_ _1843_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_8_clk_I clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5143__CLK clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4872__D Control_unit1.instr_stage1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5293__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3025__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4222__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4773__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2536__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4289__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__RN net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2864__B _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4635__I _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_2_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3820_ _1341_ _1409_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3751_ _1355_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2702_ _0559_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_199_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3682_ _1146_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2633_ _2257_ _2319_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4516__A2 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5016__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ _0514_ net264 clknet_leaf_24_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2564_ _2249_ _2238_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4303_ net29 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5283_ _0445_ net95 clknet_leaf_117_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2495_ _2145_ _2183_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4234_ _1633_ _1691_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5166__CLK clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _1601_ _1650_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5181__RN net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3116_ _0819_ _0900_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4096_ _1507_ _1596_ _1599_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_209_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4545__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3047_ _0808_ _2272_ _0851_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4204__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4998_ _0160_ net272 clknet_leaf_63_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3558__A3 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3949_ _1198_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4280__I _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__RN net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4867__D Control_unit1.instr_stage1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3191__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5172__RN net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4455__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout81 net82 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout92 net111 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5039__CLK clknet_leaf_76_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2509__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3182__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5189__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2524__A4 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout194_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3485__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5163__RN net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4910__RN net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4365__I _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4921_ _0083_ net333 clknet_leaf_40_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2996__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ _0054_ net346 clknet_leaf_44_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3803_ _1311_ _1396_ _1400_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4783_ _2084_ _0668_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_221_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2613__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3734_ _1190_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3665_ _1297_ _1289_ _1298_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2616_ _2245_ _2301_ _2291_ _2302_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3596_ _1233_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3173__A1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5335_ _0497_ net263 clknet_leaf_64_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2547_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3 _2095_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5266_ _0428_ net96 clknet_leaf_117_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2478_ _2171_ net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4217_ _1672_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5197_ _0359_ net213 clknet_leaf_83_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4673__A1 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5154__RN net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4901__RN net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4079_ _1584_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4728__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3619__I _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5331__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_238_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5393__RN net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout260 net354 net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4664__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout271 net272 net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_232_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout282 net283 net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_235_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout293 net295 net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_80_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2978__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_95_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3450_ _1141_ _1136_ _1144_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout207_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2401_ _2095_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_196_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3264__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3381_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2902__A1 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5120_ _0282_ net219 clknet_leaf_86_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_clkbuf_leaf_33_clk_I clknet_4_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5051_ _0213_ net233 clknet_leaf_71_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4655__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4002_ _1530_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_48_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4407__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__CLK clknet_leaf_110_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _0066_ net297 clknet_leaf_36_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4835_ _0037_ net284 clknet_leaf_32_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[12\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5354__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_106_clk_I clknet_4_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _0827_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3717_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _1925_ _2008_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3648_ _2143_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3579_ _1143_ _1240_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__RN net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5318_ _0480_ net261 clknet_leaf_65_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5249_ _0411_ net106 clknet_leaf_108_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5127__RN net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_10_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2518__I _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4733__I _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3385__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4871__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5227__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5118__RN net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ net18 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout157_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2881_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _1881_ _1959_ _1962_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout324_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3376__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2423__I0 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _1913_ _1903_ _1915_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3502_ _0930_ _0878_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_239_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4482_ _1774_ _1859_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3128__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3433_ _1130_ _1126_ _1131_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5357__RN net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3364_ _1006_ _1085_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _0265_ net246 clknet_leaf_79_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_174_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3295_ _1041_ _1039_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3722__I _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4628__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5109__RN net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _0196_ net237 clknet_leaf_73_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3603__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4818_ _0020_ net335 clknet_leaf_41_clk net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_222_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3367__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2414__I0 Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4749_ _0986_ _2040_ _2043_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3119__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput36 net36 Dataw_en vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput47 net47 instr_mem_addr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput58 net58 instr_mem_addr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput69 net69 write_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4875__D Control_unit1.instr_stage1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4095__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3358__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3807__I _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2711__I _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3530__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3542__I _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3080_ _2121_ _0864_ _0868_ _0877_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_212_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout274_I net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3833__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3982_ _1486_ _1523_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2933_ _0760_ _0761_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2864_ _0700_ _0701_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3349__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4603_ _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2795_ _0645_ _0648_ Stack_pointer.SP_next\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3717__I _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4010__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4534_ _0570_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2572__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4465_ _1840_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3416_ _1014_ _1117_ _1119_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4396_ _1774_ _1805_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4548__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3347_ _0977_ _1071_ _1076_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3452__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3278_ _0614_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _0179_ net238 clknet_leaf_73_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3824__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4283__I _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3588__A1 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4001__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3060__I0 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2563__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output70_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A2 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3579__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__B1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_203_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ _2261_ _2244_ _2246_ _2267_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2554__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _1699_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3201_ _2090_ _0881_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_234_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4181_ _1619_ _1656_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3132_ _2299_ _2303_ _2309_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_6390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4059__A2 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3063_ _0862_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3965_ _1465_ _1508_ _1513_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4231__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__CLK clknet_leaf_101_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2916_ _0722_ _0746_ _0749_ _0750_ _0744_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_177_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3896_ _1310_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2847_ Control_unit1.instr_stage1\[3\] _0683_ _0685_ Stack_pointer.SP\[3\] _0691_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3447__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2778_ Control_unit1.instr_stage1\[3\] _0630_ _0631_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4517_ _1887_ _1877_ _1889_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4932__CLK clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4448_ _1783_ _1841_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4379_ _1750_ _1796_ _1798_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3910__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_243_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2536__A2 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2436__I _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4213__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3750_ _1352_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout237_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2701_ _2312_ _2313_ _2329_ _2377_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3681_ _1310_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _2133_ _2282_ _2318_ _2206_ _2138_ _2272_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2527__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _0513_ net264 clknet_leaf_64_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2563_ _2251_ _2207_ _2252_ _2205_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4302_ _1306_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5282_ _0444_ net95 clknet_leaf_117_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2494_ _2160_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4098__I _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4233_ _1629_ _1690_ _1694_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_229_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ _1648_ _1649_ _1651_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3115_ _2336_ _0899_ _0902_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4095_ _1597_ _1598_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3046_ _0853_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4997_ _0159_ net272 clknet_leaf_63_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4204__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3948_ _1449_ _1496_ _1502_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3177__I _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3879_ _1358_ _1447_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3905__I _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__CLK clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__D net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5260__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4828__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4978__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3954__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_161_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__A2 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__A2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout187_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4434__A2 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4920_ _0082_ net292 clknet_leaf_38_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout354_I net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _0053_ net333 clknet_leaf_36_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4198__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3802_ _1312_ _1397_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_221_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4782_ _2170_ _0754_ _0733_ _2064_ _0709_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_207_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3945__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_7_clk_I clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3733_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3664_ _1199_ _1291_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5133__CLK clknet_leaf_87_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2615_ _2288_ _2287_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3595_ _1231_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2546_ _2204_ _2235_ _2222_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5334_ _0496_ net261 clknet_leaf_24_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2477_ _2170_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5265_ _0427_ net106 clknet_leaf_107_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5283__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4216_ _1670_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5196_ _0358_ net175 clknet_leaf_92_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4147_ _1635_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2684__A1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ _1585_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3029_ _0842_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4291__I _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5090__RN net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__D Control_unit1.instr_decoder1.A\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3164__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout250 net256 net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout261 net265 net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout272 net274 net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout283 net290 net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout294 net295 net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3370__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4416__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5006__CLK clknet_leaf_55_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5156__CLK clknet_leaf_116_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3545__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2400_ _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout102_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _1031_ _0964_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2902__A2 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5050_ _0212_ net231 clknet_leaf_71_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_211_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4655__A2 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ _1453_ _1531_ _1537_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_242_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4376__I _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3280__I _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4895__RN net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4407__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _0065_ net296 clknet_leaf_35_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4834_ _0036_ net284 clknet_leaf_32_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_72_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3918__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4765_ _2034_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3716_ _0590_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4591__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4696_ _0973_ _2006_ _2010_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3647_ _1182_ _1278_ _1283_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3578_ _1204_ _1239_ _1241_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5317_ _0479_ net263 clknet_leaf_64_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2529_ _2204_ _2146_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5248_ _0410_ net244 clknet_leaf_77_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input32_I read_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5179_ _0341_ net210 clknet_leaf_89_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5029__CLK clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5179__CLK clknet_leaf_89_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3082__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4582__A1 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5063__RN net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4637__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4196__I _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4877__RN net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2880_ net35 net46 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3376__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A1 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4550_ _1914_ _1905_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5054__RN net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2423__I1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3501_ _1182_ _1169_ _1185_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4801__RN net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3275__I _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _1770_ _1858_ _1862_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3128__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4325__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3432_ _1041_ _1128_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3363_ _0999_ _1084_ _1086_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2887__A1 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _0264_ net242 clknet_leaf_80_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3294_ _0785_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5033_ _0195_ net239 clknet_leaf_73_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2639__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__RN net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_228_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2811__A1 Stack_pointer.SP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_60_clk clknet_4_12_0_clk clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _0019_ net336 clknet_leaf_42_clk net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4564__A1 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4748_ _0801_ _2041_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4679_ _1980_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput37 net37 Serial_output vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_227_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput48 net48 instr_mem_addr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_153_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput59 net59 instr_mem_addr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2878__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_94_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4859__RN net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4744__I _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3055__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_227_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_241_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2802__A1 Stack_pointer.SP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_51_clk clknet_4_14_0_clk clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_32_clk_I clknet_4_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_47_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2869__A1 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2439__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[1\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_105_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3981_ _1480_ _1522_ _1524_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2932_ net62 _0707_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_206_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3597__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5275__RN net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_42_clk clknet_4_15_0_clk clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_241_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2863_ Arithmetic_Logic_Unit.ALU_001.p_Z _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3349__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _0966_ _1068_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2794_ Control_unit1.instr_stage1\[5\] _0630_ _0631_ _0646_ _0647_ _0648_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_157_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4533_ _1802_ _1891_ _1901_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_184_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _1838_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3415_ _1016_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3733__I _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4395_ _1770_ _1804_ _1808_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_213_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _1043_ _1073_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3277_ _1024_ _1015_ _1026_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_189_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5016_ _0178_ net198 clknet_leaf_67_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3037__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4861__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_clk clknet_4_7_0_clk clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_224_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5018__RN net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__CLK clknet_leaf_114_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3060__I1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5367__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output63_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3276__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4474__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4776__A1 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4776__B2 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__RN net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_clk clknet_4_3_0_clk clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__RN net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__I _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3200_ _0930_ _0752_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3503__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4700__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _1378_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3131_ _2312_ _2313_ _2314_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3062_ _0835_ _0587_ _0850_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4884__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4767__A1 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5248__RN net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_clk clknet_4_5_0_clk clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3964_ _1466_ _1509_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2915_ _0719_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3895_ _1459_ _1455_ _1461_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3728__I _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2846_ Control_unit2.instr_stage2\[3\] _0681_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2777_ Stack_pointer.SP\[0\] _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4516_ _1888_ _1879_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4447_ _1723_ _1839_ _1842_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3463__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4378_ _1752_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3329_ _1014_ _1062_ _1064_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_218_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4294__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4758__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3430__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3638__I _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3981__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3548__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2452__I _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _2376_ _2379_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_fanout132_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3680_ _2276_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2631_ _2317_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5350_ _0512_ net262 clknet_leaf_24_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3724__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2562_ _2165_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4301_ _1648_ _1737_ _1740_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3283__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5281_ _0443_ net106 clknet_leaf_107_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2493_ _2161_ _2163_ _2185_ _2137_ _2166_ _2135_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _1630_ _1691_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_4_clk clknet_4_4_0_clk clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ _1597_ _1650_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_229_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3114_ _0816_ _0900_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4094_ _1587_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3045_ _0805_ _2251_ _0851_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5062__CLK clknet_leaf_103_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__A2 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3660__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4996_ _0158_ net138 clknet_4_2_0_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3412__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3947_ _1501_ _1499_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_221_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3458__I _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3963__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3878_ _1293_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ _0673_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3715__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3479__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3921__I _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_226_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout83 net92 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3954__A2 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout94 net98 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2914__B1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_237_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2648__S _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3831__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout347_I net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4850_ _0052_ net335 clknet_leaf_41_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3801_ _1307_ _1396_ _1399_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4198__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4781_ _2058_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3278__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3945__A2 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3732_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3663_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2614_ _2271_ _2300_ _2286_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3594_ _1218_ _1245_ _1250_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5333_ _0495_ net271 clknet_leaf_64_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2545_ _2107_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5264_ _0426_ net251 clknet_leaf_77_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2476_ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4215_ _1606_ _1678_ _1683_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5195_ _0357_ net171 clknet_leaf_92_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4146_ _1190_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3028_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3633__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3188__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4979_ _0141_ net139 clknet_leaf_22_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_200_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3936__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3149__B1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout240 net241 net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout251 net252 net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout262 net265 net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_232_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout273 net274 net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout284 net289 net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2675__A2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout295 net301 net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4945__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3624__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3826__I _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3561__I _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4000_ _1505_ _1533_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3615__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4902_ _0064_ net299 clknet_leaf_34_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_209_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _0035_ net134 clknet_4_6_0_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_205_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5100__CLK clknet_leaf_101_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3918__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4764_ _2032_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4040__A1 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3715_ _1334_ _1335_ _1338_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4695_ _1923_ _2008_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3736__I _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5250__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3646_ _1184_ _1279_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4343__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3577_ _1138_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5316_ _0478_ net136 clknet_leaf_0_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2528_ _2175_ _2196_ _2200_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5247_ _0409_ net251 clknet_leaf_77_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2459_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[1\].i3 _2152_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5178_ _0340_ net205 clknet_leaf_94_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input25_I read_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2657__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _1623_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3909__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4889__D net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4334__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3381__I _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_clk_I clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5123__CLK clknet_leaf_116_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5273__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4799__D _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3500_ _1184_ _1172_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout212_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4480_ _1771_ _1859_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3431_ _0973_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3362_ _1001_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5101_ _0263_ net242 clknet_leaf_81_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3291__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3293_ _0962_ _1036_ _1040_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5032_ _0194_ net198 clknet_leaf_63_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2639__A2 Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2635__I _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _0018_ net334 clknet_leaf_42_clk net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4747_ _0794_ _2040_ _2042_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2575__A1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[6\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2575__B2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4678_ _1978_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3629_ _1260_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 data_mem_addr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput49 net49 instr_mem_addr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4297__I _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3827__A1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_201_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4491__A1 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2455__I _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout162_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3980_ _1482_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_223_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4243__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2931_ _0722_ _0758_ _0763_ _0750_ _0760_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_231_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_149_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2862_ Control_unit2.instr_stage2\[11\] _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4601_ _1913_ _1944_ _1949_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4546__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2793_ Stack_pointer.SP\[2\] _0642_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5019__CLK clknet_leaf_57_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4532_ _1900_ _1893_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4463_ _1747_ _1846_ _1851_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3414_ _1099_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _1771_ _1805_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3345_ _0974_ _1071_ _1075_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_217_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3276_ _1025_ _1017_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3809__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5015_ _0177_ net198 clknet_leaf_67_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2493__B1 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2493__C2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2796__A1 Stack_pointer.SP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__I _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2548__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output56_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4755__I _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3276__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4225__A1 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3200__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3130_ _2348_ _2351_ _0560_ _0563_ _2332_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_6370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__RN net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3061_ _0861_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3267__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4767__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ _1462_ _1508_ _1512_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_195_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2778__A1 Control_unit1.instr_stage1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2778__B2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2914_ _0747_ _0748_ _0727_ _2282_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_182_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3894_ _1460_ _1457_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2845_ _0689_ net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_93_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2776_ _0619_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4515_ net31 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4446_ _1779_ _1841_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4377_ _1780_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3328_ _1016_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_clk_I clknet_4_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3259_ _1011_ _1002_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_46_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4758__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2769__A1 Control_unit1.instr_stage1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4998__RN net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5334__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_104_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3194__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_119_clk_I clknet_4_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A1 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5175__RN net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4446__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3829__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3421__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4989__RN net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout125_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2630_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i0 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3185__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2561_ _2250_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3564__I _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2932__A1 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4300_ _1738_ _1739_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _0442_ net251 clknet_leaf_76_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2492_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4231_ _1626_ _1690_ _1693_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4851__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5166__RN net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4162_ _1639_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3113_ _2322_ _0899_ _0901_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4093_ _1137_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3044_ _0852_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5357__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ _0157_ net138 clknet_leaf_119_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3946_ _1195_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3877_ _1442_ _1445_ _1448_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2828_ _0625_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2759_ _0615_ net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2923__A1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4429_ _1760_ _1826_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4676__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5157__RN net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4428__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3649__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout84 net85 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout95 net97 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3384__I _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5396__RN net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2914__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2914__B2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4667__A1 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5148__RN net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3890__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3642__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ _1308_ _1397_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout242_I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4780_ net76 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_221_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3731_ _1033_ _1229_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3662_ _2188_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2613_ _2235_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3294__I _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3593_ _1166_ _1246_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5387__RN net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2905__B2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5332_ _0494_ net136 clknet_leaf_0_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2544_ _2210_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_138_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _0425_ net253 clknet_leaf_74_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2475_ _2145_ _2158_ _2168_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4214_ _1607_ _1679_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_218_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5194_ _0356_ net171 clknet_leaf_93_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4145_ _1636_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_233_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4076_ _1528_ _1286_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_243_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3027_ _0840_ _0623_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_209_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3469__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4978_ _0140_ net139 clknet_leaf_22_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4897__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3929_ _1485_ _1481_ _1487_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3149__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__RN net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout230 net259 net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout241 net258 net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_232_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3321__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout252 net253 net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout263 net265 net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout274 net279 net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout285 net288 net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout296 net298 net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3388__A1 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4003__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5052__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3312__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2458__I _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout192_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3863__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_226_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3615__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _0063_ net299 clknet_leaf_37_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3289__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _0034_ net283 clknet_leaf_32_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i0
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3379__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ _0821_ _2046_ _2051_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4040__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3714_ _1336_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_222_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4694_ _0961_ _2006_ _2009_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3645_ _1178_ _1278_ _1282_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3576_ _1233_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3551__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2527_ _2217_ _2194_ _2195_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5315_ _0477_ net130 clknet_leaf_0_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2458_ _2109_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5246_ _0408_ net243 clknet_leaf_74_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_44_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5177_ _0339_ net205 clknet_leaf_94_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2389_ Control_unit2.instr_decoder2.A\[2\] _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4128_ _1587_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input18_I read_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4059_ _1474_ _1572_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_232_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3199__I Control_unit2.instr_stage2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3927__I _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4031__A2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__CLK clknet_leaf_110_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3790__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3137__A4 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4912__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ _1123_ _1126_ _1129_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout205_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4668__I _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3533__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3361_ _1072_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5100_ _0262_ net176 clknet_leaf_101_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3292_ _1037_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ _0193_ net198 clknet_leaf_67_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3836__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4797__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4261__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4815_ _0017_ net335 clknet_leaf_42_clk net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_210_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2651__I _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _0797_ _2041_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_202_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2575__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3772__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ _1942_ _1992_ _1997_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4935__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3628_ _1258_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput39 net39 data_mem_addr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_192_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3482__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3559_ _0700_ Control_unit2.instr_stage2\[11\] _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5229_ _0391_ net214 clknet_leaf_82_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3827__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2826__I Stack_pointer.SP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4004__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3763__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3515__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3818__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4491__A2 _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5240__CLK clknet_leaf_102_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_245_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2930_ _0759_ _0748_ _0715_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout155_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2861_ Control_unit2.instr_stage2\[12\] _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout322_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4600_ _1914_ _1945_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2792_ Stack_pointer.SP\[2\] _0622_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4958__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ net20 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4462_ _1748_ _1847_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3413_ _1097_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4393_ _1767_ _1804_ _1807_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3344_ _1041_ _1073_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3275_ _0834_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _0176_ net197 clknet_leaf_66_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_227_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3285__A3 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4482__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2493__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2493__B2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4234__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3477__I _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3045__I0 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2548__A2 Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_5_clk_I clknet_4_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _0837_ _2026_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_clk clknet_4_0_0_clk clknet_leaf_110_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5113__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__I _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2757__S _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__I _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5263__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output49_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4225__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_101_clk clknet_4_9_0_clk clknet_leaf_101_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_173_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3850__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3060_ _0832_ _0566_ _0856_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2466__I _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout272_I net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2475__A1 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ _1463_ _1509_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_225_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2913_ _0712_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3297__I _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3893_ _1142_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2844_ _0688_ _0679_ _0672_ Control_unit1.instr_stage1\[2\] _0684_ Stack_pointer.SP\[2\]
+ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_176_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5136__CLK clknet_leaf_86_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2775_ _0627_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4514_ _2296_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4445_ _1840_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5286__CLK clknet_leaf_106_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4152__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4376_ _1777_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3327_ _1038_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3760__I _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3258_ _0823_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3189_ _0828_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2481__A4 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__I _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3194__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3670__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5009__CLK clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__CLK clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2560_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[6\].i3 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout118_I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2491_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[3\].i3 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4230_ _1627_ _1691_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_218_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4685__A2 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ _1636_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2696__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3112_ _0812_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4092_ _1585_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4437__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3043_ _0802_ _2273_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4994_ _0156_ net138 clknet_leaf_119_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3948__A1 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3945_ _1442_ _1496_ _1500_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3876_ _1354_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ Control_unit1.instr_stage1\[12\] Control_unit1.instr_stage1\[11\] _0674_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2758_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2923__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2689_ _2131_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[12\].i3 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4428_ _1758_ _1825_ _1829_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_232_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4586__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ net26 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4428__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_230_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout85 net88 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_161_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout96 net97 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2914__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_92_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2850__A1 Control_unit1.instr_stage1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2850__B2 Stack_pointer.SP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__RN net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3730_ _1348_ _1335_ _1350_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout235_I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2602__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_30_clk_I clknet_4_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__RN net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3661_ _1294_ _1289_ _1295_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3575__I _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _2216_ _2219_ _2298_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3592_ _1163_ _1245_ _1249_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5331_ _0493_ net131 clknet_leaf_0_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2543_ _2233_ net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_45_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5262_ _0424_ net249 clknet_leaf_74_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2474_ _2160_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _1603_ _1678_ _1682_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_218_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5193_ _0355_ net170 clknet_leaf_94_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_190_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3330__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4898__RN net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4144_ _1635_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5324__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ _1284_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_103_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3026_ net77 net78 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3094__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_90_clk clknet_4_10_0_clk clknet_leaf_90_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_180_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_118_clk_I clknet_4_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4977_ _0139_ net261 clknet_leaf_24_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5075__RN net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3928_ _1486_ _1483_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_225_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3859_ _1379_ _1430_ _1435_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout220 net221 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_236_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout231 net232 net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout242 net248 net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout253 net255 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout264 net265 net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout275 net278 net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout286 net288 net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout297 net300 net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_81_clk clknet_4_11_0_clk clknet_leaf_81_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_188_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4841__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4585__A1 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__RN net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2899__B2 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3560__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout185_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ _0062_ net287 clknet_leaf_34_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout352_I net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_72_clk clknet_4_11_0_clk clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4831_ _0033_ net148 clknet_leaf_18_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i2
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3379__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4576__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _0823_ _2047_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4804__RN net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _1290_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4693_ _1919_ _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4328__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3644_ _1180_ _1279_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3000__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3575_ _1231_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5314_ _0476_ net130 clknet_leaf_0_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2526_ _2162_ _2108_ _2104_ _2178_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3551__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout98_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5245_ _0407_ net234 clknet_leaf_71_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2457_ _2134_ _2146_ _2147_ _2150_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_229_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4500__A1 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5176_ _0338_ net159 clknet_leaf_97_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2388_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_229_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _1170_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ _1468_ _1571_ _1573_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4085__B _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4864__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2384__I Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3009_ net21 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5296__RN net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_63_clk clknet_4_12_0_clk clknet_leaf_63_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3943__I _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2559__I _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4774__I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_54_clk clknet_4_14_0_clk clknet_leaf_54_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5039__RN net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3781__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout100_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4730__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3360_ _1070_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__RN net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2469__I _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3291_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ _0192_ net197 clknet_leaf_66_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4887__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4797__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5278__RN net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_45_clk clknet_4_15_0_clk clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_207_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4814_ _0016_ net296 clknet_leaf_36_clk net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_222_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3221__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4745_ _2034_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4676_ _1900_ _1993_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3627_ _1149_ _1266_ _1271_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__RN net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3558_ Control_unit2.instr_stage2\[8\] _0752_ _0759_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2509_ _2175_ _2179_ _2200_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_5307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3489_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5228_ _0390_ net176 clknet_leaf_101_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input30_I read_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5159_ _0321_ net168 clknet_leaf_95_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5269__RN net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_clk clknet_4_13_0_clk clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3003__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5042__CLK clknet_leaf_108_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3460__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5192__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3212__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_240_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_clk clknet_4_3_0_clk clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_225_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_245_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2860_ _0698_ _0699_ net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3203__A1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2791_ Stack_pointer.SP\[2\] _0621_ _0635_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout315_I net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4530_ _1898_ _1891_ _1899_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4679__I _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ _1744_ _1846_ _1850_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3412_ _1060_ _1111_ _1116_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4703__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4392_ _1768_ _1805_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _0962_ _1071_ _1074_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3274_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2927__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _0175_ net196 clknet_leaf_66_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5065__CLK clknet_leaf_101_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18_clk clknet_4_7_0_clk clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_183_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3045__I1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2989_ net32 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4728_ _1023_ _2025_ _2029_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4589__I _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4659_ _1980_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3493__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4170__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3433__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3984__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5088__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2747__I _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout265_I net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4925__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3424__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _1459_ _1508_ _1511_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2912_ Control_unit2.instr_stage2\[8\] _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_189_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3892_ _1306_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2843_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2774_ _0626_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2935__B1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4513_ _1884_ _1877_ _1886_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_7_clk clknet_4_5_0_clk clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4444_ _1837_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4152__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4375_ _1747_ _1790_ _1795_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3326_ _1035_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3257_ _1009_ _1000_ _1010_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3188_ _0937_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3488__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4391__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4112__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__CLK clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4143__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_235_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output61_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2457__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3406__A1 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_242_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4022__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3066__C Control_unit2.instr_decoder2.A\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ _2176_ _2182_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4134__A2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3861__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4160_ _1364_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2477__I _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3111_ _0887_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _1594_ _1586_ _1595_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_237_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3042_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3645__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_4_clk_I clknet_4_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4692__I _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _0155_ net138 clknet_leaf_22_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3101__I _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3948__A2 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3944_ _1497_ _1499_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3875_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2826_ Stack_pointer.SP\[0\] _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5253__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4373__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2757_ _0611_ _0613_ _2145_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2688_ _2305_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_219_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4427_ _1800_ _1826_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_232_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4358_ _1731_ _1778_ _1784_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2687__A2 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4088__B _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3309_ _0987_ _1048_ _1051_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_219_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4289_ _1642_ _1729_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3636__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3011__I _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2611__A2 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3946__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout86 net87 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout97 net98 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_202_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__I _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3627__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5126__CLK clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5276__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2602__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2760__I Control_unit2.instr_decoder2.A\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout130_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ _1196_ _1291_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3077__B _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2611_ _2223_ _2241_ _2266_ _2287_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3591_ _1216_ _1246_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5330_ _0492_ net131 clknet_leaf_2_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2542_ _2145_ _2229_ _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4107__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5261_ _0423_ net238 clknet_leaf_73_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2473_ _2161_ _2135_ _2163_ _2164_ _2166_ _2106_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4212_ _1604_ _1679_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_218_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5192_ _0354_ net157 clknet_leaf_96_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_214_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4143_ _1528_ _1033_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4074_ _1491_ _1577_ _1582_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3025_ _0615_ _0826_ _0839_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3094__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4976_ _0138_ net344 clknet_leaf_46_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4594__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3927_ _1175_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3766__I _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3858_ _1331_ _1431_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2809_ Control_unit1.instr_stage1\[8\] _0637_ _0639_ _0658_ _0659_ _0660_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4346__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3789_ _1285_ _1389_ _1392_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout210 net216 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_236_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout221 net222 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3857__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5149__CLK clknet_leaf_87_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout232 net235 net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_232_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout243 net248 net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout254 net255 net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout265 net270 net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout276 net278 net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout287 net289 net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout298 net300 net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2845__I _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3085__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_231_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3676__I _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2755__I _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2823__A2 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4830_ _0032_ net145 clknet_leaf_17_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[7\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout345_I net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4761_ _1008_ _2046_ _2050_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2704__B _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3586__I _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2587__A1 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3712_ _1170_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4692_ _2007_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3643_ _1174_ _1278_ _1281_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3574_ _1134_ _1232_ _1238_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5313_ _0475_ net136 clknet_leaf_0_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2525_ _2120_ _2127_ _2214_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_192_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5244_ _0406_ net193 clknet_leaf_70_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2456_ _2082_ _2148_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3839__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4500__A2 _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _0337_ net157 clknet_leaf_96_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2387_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_229_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _1585_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2665__I _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _1470_ _1572_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_244_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3008_ _0778_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4959_ _0121_ net343 clknet_leaf_46_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_221_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_91_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2502__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_44_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4798__RN net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_59_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5314__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_102_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4730__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3290_ _1034_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_117_clk_I clknet_4_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout295_I net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4494__A1 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4797__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4813_ _0015_ net296 clknet_leaf_35_clk net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_222_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4744_ _2032_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4675_ _1898_ _1992_ _1996_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3626_ _1151_ _1267_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3557_ _1182_ _1220_ _1225_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2508_ _2199_ _2179_ _2181_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ net22 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _0389_ net172 clknet_leaf_93_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4831__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2439_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[1\].i3 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4485__A1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _0320_ net158 clknet_leaf_95_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input23_I read_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4109_ _1318_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5089_ _0251_ net101 clknet_leaf_109_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4981__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2799__A1 Control_unit1.instr_stage1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5337__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4115__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2723__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4785__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2790_ _0636_ _0644_ Stack_pointer.SP_next\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3203__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2962__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout210_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout308_I net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ _1745_ _1847_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3411_ _1011_ _1112_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4391_ _1762_ _1804_ _1806_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5196__RN net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3342_ _1037_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3273_ _0603_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _0174_ net186 clknet_leaf_106_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2988_ _0778_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ _0834_ _2026_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3774__I _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ _1978_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3609_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4589_ _2369_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5187__RN net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4934__RN net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3014__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3949__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4630__A1 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5111__RN net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_240_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4697__A1 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4449__A1 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout160_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3960_ _1460_ _1509_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout258_I net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4621__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__RN net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2911_ _0743_ _0745_ _0715_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2632__B1 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3891_ _1365_ _1455_ _1458_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2632__C2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2842_ _2101_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2773_ Stack_pointer.SP\[0\] _0622_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2935__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4512_ _1885_ _1879_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _1838_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5169__RN net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__CLK clknet_leaf_63_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4374_ _1748_ _1791_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2938__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3325_ _1060_ _1054_ _1061_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3256_ _0819_ _1002_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3112__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3187_ _0935_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5341__RN net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3769__I _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3415__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4612__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3179__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3009__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_239_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output54_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3103__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_246_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2457__A3 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2583__I _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5055__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4303__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3590__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3342__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2758__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3110_ _0885_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _1505_ _1588_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3041_ _0841_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3645__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4992_ _0154_ net318 clknet_leaf_54_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3943_ _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4070__A2 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3874_ _1443_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2825_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2908__A1 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2756_ _0585_ _0612_ _0601_ _2118_ _2252_ _0587_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_173_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3581__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2687_ _2364_ _2258_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4426_ _1755_ _1825_ _1828_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3333__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4357_ _1783_ _1781_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3308_ _0988_ _1049_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4288_ _1293_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3239_ _0807_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3499__I _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2844__C2 Stack_pointer.SP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2447__I0 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4061__A2 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5078__CLK clknet_leaf_102_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout76 net51 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2611__A3 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout87 net88 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout98 net110 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3572__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4915__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3324__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2578__I _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3202__I _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4033__I _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout123_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2610_ _2297_ net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3590_ _1159_ _1245_ _1248_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2541_ _2210_ _2221_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3872__I _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2472_ _2165_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5260_ _0422_ net199 clknet_leaf_67_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ _1600_ _1678_ _1681_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5191_ _0353_ net155 clknet_leaf_96_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3866__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ _1632_ _1622_ _1634_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_229_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4073_ _1492_ _1578_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3024_ _0838_ _0829_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5220__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ _0137_ net342 clknet_leaf_46_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4043__A2 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2951__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3926_ _1339_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_205_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3857_ _1329_ _1430_ _1434_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2808_ Stack_pointer.SP\[5\] _0632_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4938__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3788_ _1354_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3554__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2739_ _0595_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_195_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3306__A1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout200 net201 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4409_ _1787_ _1814_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5389_ _0551_ net322 clknet_leaf_50_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout211 net215 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout222 net229 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout233 net235 net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout244 net247 net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout255 net256 net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_232_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout266 net269 net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout277 net279 net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout288 net289 net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_235_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout299 net301 net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_189_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3085__A3 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3022__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3957__I _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_clk_I clknet_4_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3692__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4273__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4025__A2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout240_I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout338_I net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4760_ _0818_ _2047_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3711_ _1288_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4691_ _2004_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3642_ _1176_ _1279_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_220_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3573_ _1202_ _1234_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2744__C1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5312_ _0474_ net317 clknet_leaf_53_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2524_ _2105_ _2112_ _2194_ _2196_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_143_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2455_ _2098_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5243_ _0405_ net194 clknet_leaf_70_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3839__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2386_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5174_ _0336_ net155 clknet_leaf_96_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ _1333_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4056_ _1559_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4264__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3007_ _0822_ _0810_ _0825_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4016__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _0120_ net343 clknet_leaf_46_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3909_ _1468_ _1469_ _1472_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ net16 net115 clknet_leaf_6_clk Control_unit1.instr_stage1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_197_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3527__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5116__CLK clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5266__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4255__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3687__I _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2591__I _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_230_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3518__A1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4311__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4494__A2 _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout190_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout288_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4246__A2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4812_ _0014_ net299 clknet_leaf_35_clk net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_222_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4743_ _0979_ _2033_ _2039_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5139__CLK clknet_leaf_116_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4674_ _1940_ _1993_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3625_ _1145_ _1266_ _1270_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_200_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4182__A1 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5289__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3556_ _1184_ _1221_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2507_ _2134_ _2173_ _2104_ _2150_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3487_ _1019_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5226_ _0388_ net170 clknet_leaf_94_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2438_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4485__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5157_ _0319_ net174 clknet_leaf_100_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4108_ _1606_ _1596_ _1608_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_245_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5088_ _0250_ net245 clknet_leaf_78_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input16_I instr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _1501_ _1560_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3300__I _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_166_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_113_clk clknet_4_0_0_clk clknet_leaf_113_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4131__I _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4476__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4228__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4306__I _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3039__I0 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3210__I _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_104_clk clknet_4_9_0_clk clknet_leaf_104_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3410_ _1009_ _1111_ _1115_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4164__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout203_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4390_ _1764_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2714__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3341_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3272_ _1020_ _1015_ _1022_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I instr[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _0173_ net109 clknet_leaf_107_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4219__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_90_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4216__I _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3120__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ _2297_ _0796_ _0809_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4726_ _1019_ _2025_ _2028_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ _1875_ _1979_ _1985_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_200_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4155__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3608_ _1257_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4588_ _1898_ _1936_ _1941_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3539_ _1161_ _1212_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_43_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _0371_ net170 clknet_leaf_94_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_58_clk_I clknet_4_12_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5304__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_101_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4126__I _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3030__I _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_116_clk_I clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_240_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4449__A2 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3205__I _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2880__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4036__I _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2910_ _0737_ _0738_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout153_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2632__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2632__B2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ _1456_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2841_ _0682_ _0686_ net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3875__I _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4821__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout320_I net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2772_ _0626_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_223_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2935__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4511_ net30 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4442_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4971__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4688__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4373_ _1744_ _1790_ _1794_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3324_ _1011_ _1055_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5327__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3255_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3186_ _0822_ _0949_ _0954_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__A2 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2623__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3785__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4709_ _0807_ _2014_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4300__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output47_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4844__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5096__RN net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2614__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4994__CLK clknet_leaf_119_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5020__RN net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3040_ _0849_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2774__I _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout270_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2853__A1 Control_unit1.instr_stage1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2853__B2 Stack_pointer.SP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ _0153_ net317 clknet_leaf_54_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_224_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3942_ _1494_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4834__RN net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3873_ _1444_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4358__A1 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2824_ Control_unit1.instr_decoder1.A\[0\] _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2755_ _0600_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2686_ _2369_ net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2949__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _1756_ _1826_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3333__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5011__RN net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4356_ net25 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3307_ _1047_ _1048_ _1050_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4287_ _1723_ _1727_ _1730_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_189_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3238_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4867__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2844__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3169_ _0798_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2844__B2 Control_unit1.instr_stage1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_93_clk clknet_4_8_0_clk clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4597__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4825__RN net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout77 Control_unit1.instr_decoder1.A\[2\] net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2611__A4 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout88 net91 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout99 net103 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3021__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2594__I _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_84_clk clknet_4_10_0_clk clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5069__RN net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4816__RN net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3260__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3012__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5172__CLK clknet_leaf_113_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout116_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2540_ _2230_ _2164_ _2166_ _2185_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4760__A1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2471_ _2125_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ _1601_ _1679_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4512__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ _0352_ net155 clknet_leaf_96_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ _1633_ _1624_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_229_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3079__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4072_ _1488_ _1577_ _1581_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3023_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_75_clk clknet_4_14_0_clk clknet_leaf_75_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_209_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4579__A1 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ _0136_ net340 clknet_leaf_46_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4807__RN net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3925_ _1480_ _1481_ _1484_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _1376_ _1431_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2807_ Stack_pointer.SP\[5\] _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3787_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4751__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3554__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2738_ _0586_ _2259_ _0593_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5232__RN net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2669_ _2353_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ _1733_ _1812_ _1817_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5388_ _0550_ net329 clknet_leaf_29_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout201 net202 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout212 net215 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout223 net228 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout234 net235 net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4339_ _1767_ _1763_ _1769_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout245 net247 net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout256 net257 net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout267 net269 net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout278 net279 net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout289 net290 net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2817__A1 Control_unit1.instr_stage1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3303__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5045__CLK clknet_leaf_102_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_66_clk clknet_4_9_0_clk clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5195__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3793__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5223__RN net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2808__A1 Stack_pointer.SP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_57_clk clknet_4_14_0_clk clknet_leaf_57_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_219_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__D _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout233_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3710_ _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _2005_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3641_ _1168_ _1278_ _1280_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3572_ _1132_ _1232_ _1237_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2744__B1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5311_ _0473_ net317 clknet_leaf_53_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2744__C2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2523_ _2151_ _2154_ _2179_ _2181_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5242_ _0404_ net193 clknet_leaf_69_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2454_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[1\].i3 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5173_ _0335_ net163 clknet_leaf_99_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2385_ Arithmetic_Logic_Unit.ALU_000.ALU_func\[1\] _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5068__CLK clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ _1520_ _1610_ _1620_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_217_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 Serial_input net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4055_ _1557_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_48_clk clknet_4_15_0_clk clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3006_ _0824_ _0813_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3472__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4905__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4957_ _0119_ net341 clknet_leaf_48_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3908_ _1470_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3775__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ net15 net114 clknet_leaf_7_clk Control_unit1.instr_stage1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_193_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3839_ _1300_ _1417_ _1423_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2911__B _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4724__A1 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_39_clk clknet_4_13_0_clk clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2872__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4191__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5210__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_9_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout183_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4928__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3454__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3878__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2782__I _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout350_I net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _0013_ net297 clknet_leaf_36_clk net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4742_ _0791_ _2035_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_241_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4673_ _1895_ _1992_ _1995_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4502__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3624_ _1147_ _1267_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3555_ _1178_ _1220_ _1224_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4182__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ _2128_ _2172_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3486_ _1168_ _1169_ _1173_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2957__I _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5225_ _0387_ net171 clknet_leaf_94_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2437_ _2131_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5156_ _0318_ net87 clknet_leaf_116_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4107_ _1607_ _1598_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5087_ _0249_ net245 clknet_leaf_78_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_186_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _1442_ _1558_ _1561_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3445__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_2_clk_I clknet_4_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2420__A2 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4412__I _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5233__CLK clknet_leaf_108_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4173__A2 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3028__I _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5383__CLK clknet_leaf_28_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2487__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3436__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3698__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3987__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_245_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3039__I1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4164__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3340_ _1069_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3271_ _1021_ _1017_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _0172_ net108 clknet_leaf_107_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5106__CLK clknet_leaf_114_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2986_ _0808_ _0799_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4725_ _0831_ _2026_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_202_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ _1927_ _1981_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3607_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4155__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4587_ _1940_ _1937_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3538_ _1153_ _1211_ _1213_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3902__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3469_ net33 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5208_ _0370_ net163 clknet_leaf_97_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ _0301_ net85 clknet_leaf_116_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3418__A1 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4091__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_240_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5129__CLK clknet_leaf_87_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3409__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2880__A2 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4317__I _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5279__CLK clknet_leaf_76_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2632__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2840_ Control_unit1.instr_stage1\[1\] _0683_ _0685_ Stack_pointer.SP\[1\] _0686_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout146_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2771_ net77 net78 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4510_ _2276_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout313_I net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4137__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _0931_ _0966_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_208_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4372_ _1745_ _1791_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2943__I0 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3323_ _0821_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3254_ _2353_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_234_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3185_ _0824_ _0950_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2456__B _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4227__I _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2970__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2969_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4708_ _0990_ _2013_ _2017_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4639_ _1908_ _1972_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3041__I _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4064__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2614__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout263_I net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4990_ _0152_ net318 clknet_leaf_55_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3941_ _1190_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2605__A2 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_42_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3872_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2823_ _0669_ net78 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2754_ _0607_ _0608_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_57_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2685_ _2160_ _2363_ _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4510__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_100_clk_I clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4424_ _1750_ _1825_ _1827_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4355_ _1723_ _1778_ _1782_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2541__A1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3306_ _0983_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _1638_ _1729_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_115_clk_I clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2965__I _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3237_ _2296_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3097__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3062__S _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3168_ _0937_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3099_ _2213_ _0886_ _0892_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4597__A2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3796__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout78 Control_unit1.instr_decoder1.A\[1\] net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout89 net91 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_206_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3021__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4811__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__CLK clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__CLK clknet_leaf_64_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4760__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4330__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ _2136_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout109_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A2 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2523__A1 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ _1183_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4071_ _1489_ _1578_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3022_ net24 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _0135_ net340 clknet_leaf_47_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3924_ _1482_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3855_ _1325_ _1430_ _1433_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2806_ _0619_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4200__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3786_ _1387_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2737_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_199_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4240__I _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2668_ _2341_ _2352_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4407_ _1785_ _1814_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ _0549_ net329 clknet_leaf_49_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2599_ _2285_ _2286_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xfanout202 net203 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout213 net215 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout224 net228 net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_236_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout235 net241 net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4338_ _1768_ _1765_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout246 net248 net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout257 net258 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout268 net270 net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout279 net280 net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4269_ _1697_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4267__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_228_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4984__CLK clknet_leaf_63_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4019__A1 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3490__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2753__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2753__B2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4982__RN net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2505__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2808__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_5_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2992__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3640_ _1171_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout226_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3571_ _1199_ _1234_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2522_ _2213_ net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5310_ _0472_ net316 clknet_leaf_56_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2453_ _2103_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ _0403_ net231 clknet_leaf_70_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_216_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4497__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5172_ _0334_ net84 clknet_leaf_113_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_155_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2384_ Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\] _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_151_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4123_ _1619_ _1612_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3404__I _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 instr[0] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4054_ _1465_ _1565_ _1570_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_237_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3005_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5150__RN net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4956_ _0118_ net330 clknet_leaf_49_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3907_ _1446_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4887_ net14 net112 clknet_leaf_7_clk Control_unit1.instr_stage1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3838_ _1362_ _1419_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_197_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4724__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3769_ _2369_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2735__B2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5012__CLK clknet_leaf_106_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3160__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3314__I _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5162__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5141__RN net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4145__I _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2974__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3224__I _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__RN net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout176_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__A1 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4055__I _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4810_ _0012_ net286 clknet_leaf_34_clk net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout343_I net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ _0976_ _2033_ _2038_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _1896_ _1993_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3623_ _1141_ _1266_ _1269_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5199__RN net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5035__CLK clknet_leaf_57_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3554_ _1180_ _1221_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_227_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3390__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2505_ _2194_ _2196_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_239_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3485_ _1171_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2436_ _2130_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5224_ _0386_ net157 clknet_leaf_97_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout89_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__CLK clknet_leaf_113_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ _0317_ net86 clknet_leaf_116_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5371__RN net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4106_ _1150_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5086_ _0248_ net243 clknet_leaf_78_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2973__I _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4037_ _1497_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5123__RN net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4939_ _0101_ net330 clknet_leaf_49_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_205_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2708__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4937__RN net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5362__RN net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3979__I _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4633__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5058__CLK clknet_leaf_110_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3219__I _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3270_ _0831_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3124__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout293_I net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5353__RN net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3889__I _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4624__A1 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2985_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4724_ _1013_ _2025_ _2027_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4655_ _1873_ _1979_ _1984_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3606_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ net19 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3363__A1 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2968__I _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3537_ _1156_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3468_ _1004_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3115__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _0369_ net159 clknet_leaf_97_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2419_ Control_unit1.instr_decoder1.A\[0\] _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3399_ _0992_ _1106_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5344__RN net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5138_ _0300_ net84 clknet_leaf_116_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input21_I read_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_13_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5069_ _0231_ net242 clknet_leaf_81_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3418__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5200__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5350__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4918__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3106__A1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3657__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4333__I _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2770_ Control_unit1.instr_stage1\[12\] Control_unit1.instr_stage1\[11\] _0625_ _0626_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_fanout139_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3593__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout306_I net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4440_ _1773_ _1831_ _1836_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3345__A1 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_1_clk_I clknet_4_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _1741_ _1790_ _1793_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3322_ _1009_ _1054_ _1059_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3253_ _1005_ _1000_ _1007_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_224_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5326__RN net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3184_ _2354_ _0949_ _0953_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5223__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4073__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3820__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5373__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2968_ _2233_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3584__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4707_ _0804_ _2014_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_202_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2899_ Control_unit2.instr_stage2\[6\] _0713_ _0707_ _2251_ _0735_ _0736_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4638_ _1902_ _1971_ _1973_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3336__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4569_ _2233_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3992__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2401__I _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5246__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3232__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout256_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__A3 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3871_ _0879_ _1414_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2822_ net77 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2753_ _0600_ _2371_ _0609_ _2373_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2684_ _2210_ _2367_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4423_ _1752_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3869__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4354_ _1779_ _1781_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ _1038_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4285_ _1728_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3236_ _0991_ _0982_ _0993_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_246_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4238__I _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3167_ _0935_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3098_ _0792_ _0888_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2981__I _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout79 net55 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3557__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5119__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4701__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2517__C1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__CLK clknet_leaf_106_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output52_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4148__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_219_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_206_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A2 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2891__I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2756__C1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2771__A2 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3227__I _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_1_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2523__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4070_ _1485_ _1577_ _1580_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_209_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4276__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3021_ _0604_ _0826_ _0836_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3897__I _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ _0134_ net312 clknet_leaf_50_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_240_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3923_ _1446_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3854_ _1326_ _1431_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3539__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2805_ _0653_ _0656_ Stack_pointer.SP_next\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3785_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4200__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__I _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2736_ _0586_ _2259_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_246_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2667_ _2348_ _2351_ _2279_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4406_ _1731_ _1812_ _1816_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_236_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5386_ _0548_ net310 clknet_leaf_49_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2598_ _2271_ _2110_ _2280_ _2099_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_236_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout203 net204 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2976__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout214 net215 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4337_ net22 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout225 net226 net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout236 net240 net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout247 net248 net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout258 net259 net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout269 net270 net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4268_ _1661_ _1711_ _1716_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4267__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3219_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4199_ _1583_ _1671_ _1674_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2925__B _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4019__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__CLK clknet_leaf_110_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2753__A2 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3950__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__A2 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_41_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4258__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_56_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4606__I _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4430__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_114_clk_I clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2729__C1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout121_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4341__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3570_ _1130_ _1232_ _1236_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2744__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _0402_ net183 clknet_leaf_102_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2452_ _2095_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A2 _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _0333_ net80 clknet_leaf_113_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2383_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_190_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _1165_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4053_ _1466_ _1566_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput3 instr[10] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3004_ net20 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _0117_ net331 clknet_leaf_48_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_178_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ _1155_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2432__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4886_ net13 net113 clknet_leaf_7_clk Control_unit1.instr_stage1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_220_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3837_ _1297_ _1417_ _1422_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_197_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3768_ _1329_ _1372_ _1377_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2735__A2 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2719_ _0565_ _2300_ _0575_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3699_ _1160_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4951__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2499__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5369_ _0531_ net312 clknet_leaf_50_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3160__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5307__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2671__A1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_clk clknet_4_0_0_clk clknet_leaf_116_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__I _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4479__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3505__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3151__A2 Control_unit2.instr_stage2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4651__A2 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4336__I _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout169_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ _0788_ _2035_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_107_clk clknet_4_1_0_clk clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _1890_ _1992_ _1994_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3622_ _1143_ _1267_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4974__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2717__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3553_ _1174_ _1220_ _1223_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2504_ _2195_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_196_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3484_ _1127_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ _0385_ net156 clknet_leaf_96_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2435_ _2102_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ _0316_ net86 clknet_leaf_115_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4105_ _1314_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5085_ _0247_ net243 clknet_leaf_81_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_211_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4036_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2475__B _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3150__I Control_unit2.instr_stage2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4938_ _0100_ net331 clknet_leaf_40_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2405__A1 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2922__C _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4869_ Control_unit1.instr_stage1\[4\] net123 clknet_leaf_10_clk Control_unit2.instr_stage2\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4158__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2708__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2892__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4873__RN net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__CLK clknet_leaf_63_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_197_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2404__I _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3372__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3124__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout286_I net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4066__I _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__RN net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_245_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5002__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2984_ net31 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4723_ _0827_ _2026_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_241_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4654_ _1925_ _1981_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3605_ _0931_ _1229_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5152__CLK clknet_leaf_86_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4585_ _1895_ _1936_ _1939_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3536_ _1192_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5041__RN net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ _1153_ _1154_ _1158_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5206_ _0368_ net156 clknet_leaf_97_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2418_ _2105_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3398_ _0987_ _1105_ _1108_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2984__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5137_ _0299_ net90 clknet_leaf_115_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5068_ _0230_ net175 clknet_leaf_91_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input14_I instr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ _1476_ _1544_ _1548_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_244_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4855__RN net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5280__RN net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2894__I _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2617__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__CLK clknet_leaf_106_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5175__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5271__RN net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout201_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3345__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5023__RN net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _1742_ _1791_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3321_ _1058_ _1055_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3252_ _1006_ _1002_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input6_I instr[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3183_ _0819_ _0950_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2856__A1 Control_unit1.instr_stage1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2856__B2 Stack_pointer.SP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2608__A1 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4524__I _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3033__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2967_ _2213_ _0779_ _0793_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_241_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4781__A1 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _0986_ _2013_ _2016_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5262__RN net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2898_ _0733_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4637_ _1904_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3336__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4568_ _1875_ _1918_ _1928_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3519_ _1132_ _1189_ _1200_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1787_ _1869_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2847__A1 Control_unit1.instr_stage1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_96_clk clknet_4_8_0_clk clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5048__CLK clknet_leaf_102_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2847__B2 Stack_pointer.SP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4828__RN net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3272__A1 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2663__B _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5198__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3024__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4772__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__RN net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5005__RN net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3513__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_87_clk clknet_4_10_0_clk clknet_leaf_87_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_5473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4344__I _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout151_I net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _1284_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout249_I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2821_ _2086_ _0668_ _0616_ net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_220_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4763__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2752_ _2132_ _0600_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5244__RN net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_clk clknet_4_5_0_clk clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_185_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2683_ _2365_ _2137_ _2138_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3 _2366_ _2367_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4422_ _1813_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4353_ _1780_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3304_ _1035_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4284_ _1725_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3235_ _0992_ _0984_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4519__I _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3423__I _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_78_clk clknet_4_11_0_clk clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ _2213_ _0936_ _0942_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5340__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3097_ _2190_ _0886_ _0891_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2483__B _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3006__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3999_ _1451_ _1531_ _1536_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_202_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3557__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5235__RN net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2517__B1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_69_clk clknet_4_9_0_clk clknet_leaf_69_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_219_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output45_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_0_clk_I clknet_4_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_224_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_224_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2756__C2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3508__I _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5213__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2523__A3 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3720__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5363__CLK clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3243__I _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout199_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3020_ _0835_ _0829_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_clk clknet_4_2_0_clk clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3236__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4971_ _0133_ net330 clknet_leaf_49_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_240_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3922_ _1170_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3853_ _1319_ _1430_ _1432_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2804_ Control_unit1.instr_stage1\[7\] _0630_ _0631_ _0654_ _0655_ _0656_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4736__A1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5217__RN net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2735_ _0586_ _2371_ _0592_ _2373_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2666_ _2349_ _2350_ _2343_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _1783_ _1814_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5385_ _0547_ net329 clknet_leaf_39_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2597_ _2271_ _2146_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout204 net260 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4336_ _1339_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout215 net216 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout226 net228 net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_236_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout237 net240 net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4249__I _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout248 net257 net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3153__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout259 net260 net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4267_ _1619_ _1712_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3218_ _2212_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3475__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4198_ _1638_ _1673_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3149_ _0702_ _0864_ _0920_ _0929_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_215_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3778__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4712__I _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5208__RN net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3466__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4718__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2729__B1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2729__C2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3238__I _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout114_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2520_ _2211_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2451_ _2141_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5170_ _0332_ net83 clknet_leaf_113_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2382_ Arithmetic_Logic_Unit.ALU_000.ALU_func\[0\] _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4121_ _1617_ _1610_ _1618_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4052_ _1462_ _1565_ _1569_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 instr[11] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3003_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3209__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4954_ _0116_ net337 clknet_leaf_40_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5259__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3905_ _1444_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ net12 net112 clknet_leaf_7_clk Control_unit1.instr_stage1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4709__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3836_ _1360_ _1419_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4185__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3767_ _1376_ _1373_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_238_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2718_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3932__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3698_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2649_ _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5368_ _0530_ net275 clknet_leaf_61_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2499__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3696__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4319_ _1750_ _1751_ _1754_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5299_ _0461_ net130 clknet_leaf_1_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2428__S _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3999__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2655__C _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2671__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3620__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4176__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3151__A3 Control_unit2.instr_stage2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3439__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3521__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2662__A2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3611__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout231_I net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _1892_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout329_I net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3621_ _1204_ _1266_ _1268_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4167__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3552_ _1176_ _1221_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2503_ _2184_ _2107_ _2147_ _2193_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3483_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _0384_ net155 clknet_leaf_97_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2434_ _2113_ _2128_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5153_ _0315_ net161 clknet_leaf_98_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_155_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4104_ _1603_ _1596_ _1605_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5084_ _0246_ net213 clknet_leaf_82_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4035_ _1556_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3431__I _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5081__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ _0099_ net330 clknet_leaf_40_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3602__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_40_clk_I clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4868_ Control_unit1.instr_stage1\[3\] net124 clknet_leaf_9_clk Control_unit2.instr_stage2\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4158__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3819_ _1334_ _1408_ _1410_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4799_ _0001_ net118 clknet_leaf_6_clk net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_55_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3669__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_113_clk_I clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3341__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4397__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_231_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4172__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4149__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3516__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout181_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3251__I _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout279_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3832__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4941__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2983_ _2277_ _0796_ _0806_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _2007_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4653_ _1871_ _1979_ _1983_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3604_ _1182_ _1251_ _1256_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_200_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4584_ _1896_ _1937_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3535_ _1188_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3426__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3466_ _1156_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout94_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2417_ _2106_ _2108_ _2100_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5205_ _0367_ net164 clknet_leaf_99_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3397_ _0988_ _1106_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_233_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5136_ _0298_ net219 clknet_leaf_86_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5067_ _0229_ net211 clknet_leaf_91_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_211_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4018_ _1518_ _1545_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4551__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output75_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4814__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4964__CLK clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2617__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3814__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2415__I _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3246__I _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3320_ _0818_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3251_ _0815_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3182_ _2336_ _0949_ _0952_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4077__I _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_227_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2608__A2 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3281__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2966_ _0792_ _0783_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4705_ _0801_ _2014_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2897_ net56 _0724_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2792__A1 Stack_pointer.SP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__I _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4636_ _1953_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4837__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3156__I _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _1927_ _1921_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3518_ _1199_ _1193_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _2212_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2995__I _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3449_ _1143_ _1139_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_213_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4987__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ _0281_ net220 clknet_leaf_85_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3272__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4772__A2 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2535__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__CLK clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__I _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout144_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2820_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5292__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2751_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[0\].i2 _2260_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_223_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout311_I net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2682_ _2356_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_195_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _1811_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2526__A1 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4352_ _1776_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_236_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3303_ _0794_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4283_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3234_ _0804_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_234_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3165_ _0792_ _0938_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__RN net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3096_ _0789_ _0888_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_208_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4535__I _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__C _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4451__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3998_ _1503_ _1533_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2949_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4270__I _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4994__RN net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4619_ _1882_ _1960_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2517__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2517__B2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5015__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5165__CLK clknet_leaf_87_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5171__RN net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4445__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4180__I _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2756__B2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3181__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3524__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4681__A1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout261_I net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4970_ _0132_ net337 clknet_leaf_40_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3921_ _1444_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2444__B1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2444__C2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3852_ _1321_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_242_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2803_ Stack_pointer.SP\[4\] _0632_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_220_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3783_ _0879_ _0966_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2734_ _2132_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[14\].i3 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4976__RN net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2665_ _2347_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4404_ _1723_ _1812_ _1815_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2596_ _2280_ _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5384_ _0546_ net276 clknet_leaf_29_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_246_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5188__CLK clknet_leaf_113_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout205 net210 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4335_ _1762_ _1763_ _1766_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3434__I _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout216 net230 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout227 net228 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout238 net240 net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout249 net256 net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4266_ _1617_ _1711_ _1715_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3217_ _0977_ _0969_ _0978_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5153__RN net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3148_ _0865_ _0611_ _0864_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_216_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ _0865_ _0875_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2986__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4727__A2 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3609__I _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3163__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3466__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2729__B2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2450_ _2144_ net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout107_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3154__A1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3254__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ _1518_ _1612_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4051_ _1463_ _1566_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4654__A1 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 instr[12] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_237_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3002_ _2369_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A1 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ _0115_ net337 clknet_leaf_40_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_196_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ _1318_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4884_ net11 net114 clknet_leaf_7_clk Control_unit1.instr_stage1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_221_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3835_ _1294_ _1417_ _1421_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3766_ _1215_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2717_ _0565_ _2300_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3697_ _2334_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2648_ _2332_ _2333_ _2141_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3145__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5367_ _0529_ net275 clknet_leaf_61_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2579_ _2261_ _2244_ _2246_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5374__RN net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4318_ _1752_ _1753_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5298_ _0460_ net130 clknet_leaf_1_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_5_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4249_ _1697_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__RN net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5203__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2959__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__D Control_unit1.instr_stage1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_204_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5353__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3339__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5117__RN net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2647__B1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2647__C2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3611__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3249__I _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout224_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3620_ _1138_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3375__A1 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3551_ _1168_ _1220_ _1222_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2502_ _2184_ _2173_ _2191_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3482_ net21 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3127__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5221_ _0383_ net162 clknet_leaf_99_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2433_ _2120_ _2127_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4870__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5152_ _0314_ net219 clknet_leaf_86_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ _1604_ _1598_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5083_ _0245_ net212 clknet_leaf_82_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3712__I _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A1 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5226__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4034_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4936_ _0098_ net293 clknet_leaf_29_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3602__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ Control_unit1.instr_stage1\[2\] net143 clknet_leaf_17_clk Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3818_ _1336_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4798_ _0000_ net119 clknet_leaf_11_clk net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_197_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3366__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2998__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3749_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3118__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3669__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4865__D Control_unit1.instr_stage1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4618__A1 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3357__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4893__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5249__CLK clknet_leaf_108_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4609__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout174_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3832__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout341_I net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2982_ _0805_ _0799_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_226_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ _2005_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ _1923_ _1981_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3348__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 read_data[6] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3603_ _1184_ _1252_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4583_ _1890_ _1936_ _1938_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3899__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3534_ _1149_ _1205_ _1210_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3465_ _1127_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5204_ _0366_ net93 clknet_leaf_110_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2416_ _2092_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout87_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3396_ _1047_ _1105_ _1107_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5135_ _0297_ net220 clknet_leaf_86_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3442__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5066_ _0228_ net232 clknet_leaf_70_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4076__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4017_ _1473_ _1544_ _1547_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3823__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_240_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3587__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4919_ _0081_ net292 clknet_leaf_37_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_209_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2521__I _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output68_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3511__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_236_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4067__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4183__I _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3578__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3250_ _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2587__B _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout291_I net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3181_ _0816_ _0950_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3262__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3805__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_54_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4093__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_223_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3569__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2965_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4230__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4704_ _1929_ _2013_ _2015_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_202_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_69_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2896_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4635_ _1951_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_112_clk_I clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3437__I _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4566_ net27 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3517_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _1873_ _1867_ _1874_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_235_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3448_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _1028_ _1090_ _1095_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _0280_ net225 clknet_leaf_85_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_246_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5049_ _0211_ net233 clknet_leaf_82_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3900__I _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5094__CLK clknet_leaf_103_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2535__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2426__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2870__B net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2750_ _0583_ _0595_ _0605_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA_fanout137_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2681_ _2364_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_195_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout304_I net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _1747_ _1819_ _1824_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2526__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4351_ net18 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3302_ _0980_ _1036_ _1046_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4282_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3233_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3164_ _2190_ _0936_ _0941_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3095_ _2171_ _0886_ _0890_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_242_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A2 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3997_ _1449_ _1531_ _1535_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4203__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2948_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3167__I _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2879_ Control_unit2.instr_stage2\[4\] _0713_ _0715_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_159_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _1929_ _1959_ _1961_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4954__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2517__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4549_ net24 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3190__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4873__D Control_unit1.instr_stage1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2447__S _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2756__A2 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2508__A2 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3705__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__A2 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__I _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4827__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4433__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout254_I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3920_ _1333_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2444__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2444__B2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ _1418_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2802_ Stack_pointer.SP\[4\] _0642_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3782_ _1348_ _1381_ _1386_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4977__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2733_ _0591_ net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2664_ _2299_ _2303_ _2309_ _2327_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_146_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4403_ _1779_ _1814_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5383_ _0545_ net276 clknet_leaf_28_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2595_ _2282_ _2164_ _2166_ _2250_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_236_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4334_ _1764_ _1765_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout206 net209 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout217 net218 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout228 net229 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4265_ _1659_ _1712_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout239 net240 net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3216_ _0789_ _0971_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4196_ _1669_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3147_ _0585_ _0702_ _0927_ _2234_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2683__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2683__B2 Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3078_ _0688_ _0871_ _0874_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4424__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2738__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4868__D Control_unit1.instr_stage1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5132__CLK clknet_leaf_90_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4360__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output50_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2685__B _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3360__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_119_clk clknet_4_2_0_clk clknet_leaf_119_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2729__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3535__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4050_ _1459_ _1565_ _1568_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3001_ _2354_ _0810_ _0820_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_232_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4366__I _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 instr[13] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3270__I _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__RN net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4406__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ _0114_ net294 clknet_leaf_38_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2417__A1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__CLK clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3903_ _1465_ _1455_ _1467_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4883_ net10 net112 clknet_leaf_7_clk Control_unit1.instr_stage1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3834_ _1358_ _1419_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__CLK clknet_leaf_116_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3765_ _1325_ _1372_ _1375_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_203_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ _0565_ _2371_ _0574_ _2373_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4590__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3696_ _1319_ _1320_ _1323_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2647_ _2133_ _2318_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3 _2206_ _2165_ _2281_
+ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3145__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5366_ _0528_ net277 clknet_leaf_28_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2578_ _2266_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4317_ _1728_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5297_ _0459_ net104 clknet_leaf_118_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_64_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4248_ _1594_ _1698_ _1704_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4645__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2656__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4179_ _1617_ _1655_ _1660_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_216_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3081__A1 Control_unit2.instr_stage2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2895__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3090__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2647__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2647__B2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5028__CLK clknet_leaf_106_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4876__RN net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5178__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3375__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4572__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3550_ _1171_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_196_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2501_ _2082_ _2192_ _2098_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4800__RN net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3265__I _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3481_ _1125_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3127__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _0382_ net81 clknet_leaf_112_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_157_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2432_ _2079_ _2123_ _2126_ _2080_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5151_ _0313_ net220 clknet_leaf_85_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2886__A1 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4102_ _1146_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5082_ _0244_ net233 clknet_leaf_82_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2609__I _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4867__RN net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4935_ _0097_ net276 clknet_leaf_29_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ Control_unit1.instr_stage1\[1\] net146 clknet_leaf_14_clk Arithmetic_Logic_Unit.ALU_000.ALU_func\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_221_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3817_ _1390_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4797_ _0710_ _2074_ _2077_ _0750_ _2075_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_222_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3748_ _2233_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ _1307_ _1302_ _1309_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_238_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5349_ _0511_ net264 clknet_leaf_25_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2877__A1 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4881__D net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5320__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3054__A1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__A1 Stack_pointer.SP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_50_clk clknet_4_13_0_clk clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4849__RN net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3293__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout167_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2981_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout334_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__A1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4720_ _1942_ _2019_ _2024_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_203_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__RN net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_clk clknet_4_15_0_clk clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_203_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4651_ _1864_ _1979_ _1982_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput20 read_data[11] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3602_ _1178_ _1251_ _1255_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput31 read_data[7] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_204_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4582_ _1892_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3533_ _1151_ _1206_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5203_ _0365_ net93 clknet_leaf_112_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2415_ _2109_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_233_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2859__A1 Control_unit1.instr_stage1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3395_ _0983_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3723__I _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2859__B2 Stack_pointer.SP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5134_ _0296_ net225 clknet_leaf_85_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5343__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5065_ _0227_ net193 clknet_leaf_101_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _1474_ _1545_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_226_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4554__I _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_226_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _0080_ net291 clknet_leaf_37_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_32_clk clknet_4_7_0_clk clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4849_ _0051_ net334 clknet_leaf_36_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_194_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5017__RN net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4876__D Control_unit1.instr_stage1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_99_clk clknet_4_8_0_clk clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_216_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4464__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4860__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4775__A1 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5256__RN net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4527__A1 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5008__RN net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5216__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5366__CLK clknet_leaf_28_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_239_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3180_ _2322_ _0949_ _0951_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_234_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout284_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4766__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5247__RN net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2964_ net27 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_14_clk clknet_4_5_0_clk clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ _0797_ _2014_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2895_ _0618_ _0706_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3718__I _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4634_ _1942_ _1965_ _1970_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4565_ _1873_ _1918_ _1926_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3516_ net26 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3741__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4496_ _1785_ _1869_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3447_ net29 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3453__I _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3378_ _1029_ _1091_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_246_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5117_ _0279_ net217 clknet_leaf_90_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5048_ _0210_ net191 clknet_leaf_102_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3257__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I instr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4883__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4757__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5239__CLK clknet_leaf_104_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3628__I _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3980__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3496__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3248__A1 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4194__I _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3799__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4748__A1 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2680_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[12\].i3 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4350_ _1777_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2526__A3 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2931__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3301_ _1045_ _1039_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4281_ _1724_ _1186_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3273__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3232_ _2276_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_3_clk clknet_4_4_0_clk clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input4_I instr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3163_ _0789_ _0938_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_230_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3094_ _0786_ _0888_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_223_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4739__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3996_ _1501_ _1533_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_241_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_241_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2947_ _0670_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3411__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3448__I _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3962__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2878_ net54 _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4617_ _1878_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3714__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4548_ _0614_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4279__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4479_ _1767_ _1858_ _1861_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3478__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3911__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3650__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3402__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_53_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4130__A2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_68_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_111_clk_I clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2437__I _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2444__A2 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3641__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3850_ _1416_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout247_I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2801_ Stack_pointer.SP\[4\] _0622_ _0635_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_220_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3781_ _1349_ _1382_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3268__I _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2732_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2663_ _2330_ _2344_ _2347_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4402_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2594_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5382_ _0544_ net277 clknet_leaf_28_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4333_ _1728_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout207 net209 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_173_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout218 net222 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4264_ _1614_ _1711_ _1714_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout229 net230 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_214_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3215_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4121__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4195_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5084__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3146_ _2139_ _0613_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2683__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A1 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3077_ _0871_ _0874_ _0688_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_215_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3632__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4921__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3178__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3979_ _1498_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3906__I _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4884__D net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3871__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3623__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_215_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4179__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3088__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3816__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4647__I _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4103__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout197_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3000_ _0819_ _0813_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 instr[14] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4944__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _0113_ net292 clknet_leaf_37_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2417__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3614__A1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4382__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3902_ _1466_ _1457_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4882_ net9 net114 clknet_leaf_7_clk Control_unit1.instr_stage1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3833_ _1285_ _1417_ _1420_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3764_ _1326_ _1373_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2715_ _2131_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[13\].i3 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3726__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3695_ _1321_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2630__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2646_ _2310_ _2328_ _2330_ _2331_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4342__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2577_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5365_ _0527_ net277 clknet_leaf_28_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4316_ net32 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5296_ _0458_ net252 clknet_leaf_78_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4557__I _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3461__I _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4247_ _1646_ _1700_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4178_ _1659_ _1656_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3853__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3129_ _0615_ _0905_ _0910_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_228_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__A1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3081__A2 Control_unit2.instr_stage2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3908__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4817__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3371__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4967__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2647__A2 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4021__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2450__I _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2500_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[3\].i3 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3480_ _1013_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2431_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_237_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _0312_ net225 clknet_leaf_85_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4101_ _1310_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4377__I _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _0243_ net233 clknet_leaf_82_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4032_ _1528_ _0931_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2638__A2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4934_ _0096_ net291 clknet_leaf_29_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_206_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4865_ Control_unit1.instr_stage1\[0\] net146 clknet_leaf_14_clk Arithmetic_Logic_Unit.ALU_000.ALU_func\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_107_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3816_ _1388_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5272__CLK clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ Control_unit2.instr_stage2\[3\] _0748_ _0714_ _2076_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_140_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3456__I _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3747_ _1300_ _1353_ _1363_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2574__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3678_ _1308_ _1304_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2629_ _2310_ _2315_ _2279_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5348_ _0510_ net137 clknet_leaf_21_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2877__A2 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5279_ _0441_ net252 clknet_leaf_76_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_211_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2565__A1 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4197__I _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__CLK clknet_leaf_87_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4490__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2980_ net30 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5295__CLK clknet_leaf_77_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ _1919_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout327_I net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput10 instr[2] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_238_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3601_ _1180_ _1252_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput21 read_data[12] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput32 read_data[8] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4581_ _1920_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3532_ _1145_ _1205_ _1209_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_196_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3463_ net32 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5202_ _0364_ net93 clknet_leaf_112_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_237_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2414_ Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\] _2078_ _2081_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3394_ _1099_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _0295_ net217 clknet_leaf_87_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5143__D _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5064_ _0226_ net173 clknet_leaf_100_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _1468_ _1544_ _1546_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4917_ _0079_ net291 clknet_leaf_37_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4784__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4570__I _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4848_ _0050_ net298 clknet_leaf_42_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4779_ _2062_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2547__A1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5018__CLK clknet_leaf_57_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3914__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5168__CLK clknet_leaf_86_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4745__I _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4472__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4224__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2786__A1 Stack_pointer.SP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2538__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__RN net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout277_I net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3266__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2963_ _2190_ _0779_ _0790_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4766__A2 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2777__A1 Stack_pointer.SP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _2007_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2894_ _0719_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _1900_ _1966_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4564_ _1925_ _1921_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3515_ _1130_ _1189_ _1197_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5310__CLK clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4495_ _2189_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3734__I _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout92_I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3446_ _0986_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3377_ _1024_ _1090_ _1094_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5183__RN net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _0278_ net211 clknet_leaf_91_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_246_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _0209_ net191 clknet_leaf_102_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_228_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2768__A1 Control_unit1.instr_stage1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4997__RN net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3193__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2940__A1 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output73_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3496__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5174__RN net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4475__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3420__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4988__RN net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5333__CLK clknet_leaf_64_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2931__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3300_ _0791_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _0965_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3231_ _0987_ _0982_ _0989_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5165__RN net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3162_ _2171_ _0936_ _0940_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4912__RN net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4385__I _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3093_ _2144_ _0886_ _0889_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_236_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_223_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3995_ _1442_ _1531_ _1534_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _0624_ _0775_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2877_ net47 net76 net52 net53 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _1953_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3175__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4547_ _1910_ _1903_ _1912_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3464__I _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2922__A1 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2922__B2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4478_ _1768_ _1859_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3429_ _1037_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4675__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3478__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4427__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5356__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3639__I _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2543__I _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_224_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5395__RN net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3641__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3549__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2800_ _0649_ _0652_ Stack_pointer.SP_next\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout142_I net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3780_ _1344_ _1381_ _1385_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2731_ _2257_ _0584_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2662_ _2345_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_246_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _1810_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5381_ _0543_ net277 clknet_leaf_28_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3284__I Control_unit2.instr_stage2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2593_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5386__RN net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4332_ net21 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout208 net209 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout219 net221 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4263_ _1615_ _1712_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4657__A1 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__RN net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5229__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3214_ _2189_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4194_ _1669_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3145_ _0567_ _0588_ _0602_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_214_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3076_ _0872_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5310__RN net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3978_ _1495_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3396__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2929_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3148__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5377__RN net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3922__I _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3871__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3387__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2448__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3311__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput8 instr[15] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3862__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4950_ _0112_ net295 clknet_leaf_30_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3901_ _1150_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4881_ net2 net112 clknet_leaf_7_clk Control_unit1.instr_stage1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3279__I _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3832_ _1354_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3763_ _1319_ _1372_ _1374_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2714_ _2364_ _2260_ _2374_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3694_ _1290_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2645_ _2323_ _2327_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_220_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5051__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5364_ _0526_ net139 clknet_leaf_22_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2576_ _2262_ _2264_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ _1726_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3742__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5295_ _0457_ net251 clknet_leaf_77_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4246_ _1592_ _1698_ _1703_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3302__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4177_ _1215_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3128_ _0838_ _0906_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_215_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3059_ _0860_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_52_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3369__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3917__I _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4030__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_67_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__A2 Arithmetic_Logic_Unit.ALU_001.Y_CY\[7\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_110_clk_I clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4021__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5074__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2430_ _2078_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout105_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3532__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4658__I _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4100_ _1600_ _1596_ _1602_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4911__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5080_ _0242_ net191 clknet_leaf_101_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4031_ _1491_ _1550_ _1555_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_238_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3835__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_206_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4796__B1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _0095_ net276 clknet_leaf_29_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_221_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4864_ _0058_ net145 clknet_leaf_17_clk Arithmetic_Logic_Unit.ALU_001.p_Z vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3815_ _1379_ _1402_ _1407_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4795_ _2075_ _2068_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _1362_ _1356_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2574__A2 Arithmetic_Logic_Unit.ALU_001.Y_CY\[6\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3771__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3677_ _1142_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2628_ _2312_ _2313_ _2314_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_66_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3523__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5347_ _0509_ net134 clknet_leaf_2_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2559_ _2159_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2877__A3 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5278_ _0440_ net249 clknet_leaf_74_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input35_I start vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4229_ _1621_ _1690_ _1692_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4251__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5097__CLK clknet_leaf_101_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3062__I0 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4934__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3514__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3382__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4490__A2 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2726__I _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4242__A2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_203_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3600_ _1174_ _1251_ _1254_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput11 instr[3] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput22 read_data[13] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4580_ _1917_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput33 read_data[9] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3531_ _1147_ _1206_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3462_ _1125_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5201_ _0363_ net89 clknet_leaf_114_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2413_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4388__I _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3393_ _1097_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _0294_ net208 clknet_leaf_90_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5063_ _0225_ net173 clknet_leaf_100_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_238_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4014_ _1470_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_238_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4481__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2636__I _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4807__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4916_ _0078_ net282 clknet_leaf_30_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4847_ _0049_ net297 clknet_leaf_36_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_194_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _0719_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2547__A2 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3729_ _1349_ _1337_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4298__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3930__I _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2483__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_231_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_clk clknet_4_8_0_clk clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5112__CLK clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3840__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5262__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout172_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2474__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4215__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2962_ _0789_ _0783_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2777__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4701_ _2005_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A1 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2893_ net56 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3287__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2405__B _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4632_ _1898_ _1965_ _1969_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_204_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2529__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4563_ net26 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3514_ _1196_ _1193_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4494_ _1871_ _1867_ _1872_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3445_ _1047_ _1136_ _1140_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_170_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3376_ _1025_ _1091_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout85_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _0277_ net211 clknet_leaf_91_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_246_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3750__I _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5046_ _0208_ net192 clknet_leaf_102_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4581__I _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3197__I _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5135__CLK clknet_leaf_86_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5285__CLK clknet_leaf_106_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output66_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3708__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2931__A2 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3230_ _0988_ _0984_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4684__A2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3161_ _0786_ _0938_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3092_ _0781_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__A2 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5008__CLK clknet_leaf_55_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3994_ _1497_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_222_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2945_ Control_unit1.instr_stage1\[0\] _0674_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5158__CLK clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2876_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4615_ _1951_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3745__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4546_ _1911_ _1905_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ _1762_ _1858_ _1860_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4124__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3428_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3359_ _0995_ _1078_ _1083_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3480__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _0191_ net196 clknet_leaf_66_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_227_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3650__A3 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5092__RN net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3655__I _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3166__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4418__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5300__CLK clknet_leaf_119_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_204_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2730_ _2257_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout135_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__RN net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2661_ _2101_ _2136_ _2339_ _2147_ _2338_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_195_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4400_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout302_I net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4354__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ _0542_ net268 clknet_leaf_26_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2592_ _2124_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[7\].i3 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _1726_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout209 net210 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4262_ _1609_ _1711_ _1713_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_218_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4657__A2 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3213_ _0974_ _0969_ _0975_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2909__I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__A1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4193_ _0883_ _1068_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3144_ _2284_ _0923_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_228_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4409__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3075_ _0612_ _2260_ _0610_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_227_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3093__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2840__A1 Control_unit1.instr_stage1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2840__B2 Stack_pointer.SP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3977_ _1520_ _1514_ _1521_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5074__RN net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2928_ net58 net59 _0742_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_210_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2859_ Control_unit1.instr_stage1\[7\] _0672_ _0684_ Stack_pointer.SP\[7\] _0699_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4529_ _1800_ _1893_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2819__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5342__D _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5323__CLK clknet_leaf_57_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3084__A1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_80_clk clknet_4_11_0_clk clknet_leaf_80_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_187_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__RN net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4812__RN net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3139__A2 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4879__RN net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 instr[1] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_237_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3075__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3900_ _1314_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4880_ Control_unit1.instr_decoder1.A\[2\] net144 clknet_leaf_16_clk Control_unit2.instr_decoder2.A\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_71_clk clknet_4_11_0_clk clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_233_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3831_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4840__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3378__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3762_ _1321_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5056__RN net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2713_ _2379_ _0559_ _2376_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4803__RN net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3693_ _1155_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2644_ _2312_ _2313_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4990__CLK clknet_leaf_55_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _0525_ net141 clknet_leaf_21_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2575_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[6\].i3 _2152_ _2263_ _2149_ _2264_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3550__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _1318_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5294_ _0456_ net249 clknet_leaf_74_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4245_ _1644_ _1700_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4176_ _1614_ _1655_ _1658_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3127_ _0604_ _0905_ _0909_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3066__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3058_ _0828_ _2365_ _0856_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_227_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5295__RN net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2813__A1 Control_unit1.instr_stage1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_clk clknet_4_12_0_clk clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4764__I _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4863__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2804__A1 Control_unit1.instr_stage1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__RN net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_53_clk clknet_4_14_0_clk clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_128_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5038__RN net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5219__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5369__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _1492_ _1551_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_238_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3296__A1 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4796__A1 Control_unit2.instr_stage2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4932_ _0094_ net266 clknet_leaf_27_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3599__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5277__RN net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_44_clk clknet_4_15_0_clk clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_240_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4863_ Stack_pointer.SP_next\[7\] net122 clknet_leaf_11_clk Stack_pointer.SP\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3814_ _1331_ _1403_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5029__RN net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4794_ net53 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3220__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3745_ _1201_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3676_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2627_ _2304_ _2308_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_6509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4720__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5201__RN net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2558_ _2242_ _2247_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_217_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5346_ _0508_ net134 clknet_leaf_2_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2877__A4 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2489_ _2179_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5277_ _0439_ net238 clknet_leaf_72_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_173_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4228_ _1623_ _1691_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input28_I read_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ _1594_ _1637_ _1647_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4787__A1 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_35_clk clknet_4_13_0_clk clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_197_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3062__I1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3663__I _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4778__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2943__S _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5259__RN net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_clk clknet_4_3_0_clk clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5041__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3450__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5191__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput12 instr[4] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput23 read_data[14] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput34 reset net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_196_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3530_ _1141_ _1205_ _1208_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout215_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4669__I _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3461_ _0998_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2412_ _2094_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5200_ _0362_ net223 clknet_leaf_83_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3392_ _0980_ _1098_ _1104_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _0293_ net208 clknet_leaf_89_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5062_ _0224_ net182 clknet_leaf_103_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _1532_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2917__I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_66_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_198_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_17_clk clknet_4_7_0_clk clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4915_ _0077_ net282 clknet_leaf_31_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3748__I _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2652__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4846_ _0048_ net296 clknet_leaf_35_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4777_ net35 _2059_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3744__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3728_ _1183_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3483__I _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3659_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_19_clk_I clknet_4_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5329_ _0491_ net136 clknet_leaf_0_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_5616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5064__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2483__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3432__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_237_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3983__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4901__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4489__I _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3393__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_226_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout165_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2961_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout332_I net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4700_ _0979_ _2006_ _2012_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2892_ _0722_ _0726_ _0728_ _0720_ _0729_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4631_ _1940_ _1966_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ _1871_ _1918_ _1924_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3513_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4493_ _1783_ _1869_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_6_clk clknet_4_5_0_clk clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3444_ _1138_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3375_ _1020_ _1090_ _1093_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5087__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _0276_ net205 clknet_leaf_88_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_218_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5045_ _0207_ net192 clknet_leaf_102_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_211_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4924__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3965__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _0031_ net148 clknet_leaf_18_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[6\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4390__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4102__I _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3941__I _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output59_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2916__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2392__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4012__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4133__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3851__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3160_ _2144_ _0936_ _0939_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2467__I _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout282_I net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3091_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4947__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3644__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3993_ _1532_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2944_ _0769_ _0720_ _0711_ _0774_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_206_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2875_ _0667_ _0706_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4614_ _1875_ _1952_ _1958_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4545_ net23 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4476_ _1764_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3427_ _1124_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4124__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3761__I _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3358_ _0996_ _1079_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3289_ _0780_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5028_ _0190_ net186 clknet_leaf_106_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input10_I instr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4592__I _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3938__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__CLK clknet_leaf_108_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3671__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3626__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3929__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2660_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3 _2096_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout128_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_201_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2591_ _2278_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_201_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ _1333_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _1611_ _1712_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3212_ _0786_ _0971_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I instr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4192_ _1632_ _1663_ _1668_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3143_ _2319_ _2333_ _2340_ _2367_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_171_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3074_ _0583_ _0605_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3617__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5125__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3093__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4290__A1 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4042__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3976_ _1478_ _1515_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2927_ net48 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2858_ Control_unit2.instr_stage2\[7\] _0679_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2789_ Control_unit1.instr_stage1\[4\] _0638_ _0640_ _0641_ _0643_ _0644_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_219_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4528_ _2353_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4459_ _1741_ _1846_ _1849_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4281__A1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2570__I _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2595__A1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5148__CLK clknet_leaf_90_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3075__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3830_ _1415_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3761_ _1355_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3576__I _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2586__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2712_ _0571_ net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_203_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3692_ _1288_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2643_ _2309_ _2327_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5362_ _0524_ net141 clknet_leaf_21_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2574_ _2130_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[6\].i3 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4313_ _1747_ _1737_ _1749_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5293_ _0455_ net234 clknet_leaf_71_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4244_ _1590_ _1698_ _1702_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4175_ _1615_ _1656_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3126_ _0835_ _0906_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3057_ _0859_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3066__A2 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3959_ _1507_ _1508_ _1510_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4110__I _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4780__I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4309__A2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout195_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4245__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4931_ _0093_ net266 clknet_leaf_25_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4796__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4690__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4862_ Stack_pointer.SP_next\[6\] net115 clknet_leaf_8_clk Stack_pointer.SP\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_146_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3813_ _1329_ _1402_ _1406_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4793_ _2212_ _0754_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3744_ _1297_ _1353_ _1361_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5313__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3675_ _2255_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2626_ _2245_ _2301_ _2291_ _2302_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _0507_ net137 clknet_leaf_21_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _2244_ _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2731__A1 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5276_ _0438_ net199 clknet_leaf_67_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2488_ _2162_ _2173_ _2180_ _2178_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__4960__RN net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4227_ _1672_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4158_ _1646_ _1640_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3109_ _2297_ _0893_ _0898_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4089_ _1299_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4236__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__A1 Stack_pointer.SP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4539__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4105__I _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2789__A1 Control_unit1.instr_stage1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5336__CLK clknet_leaf_64_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_8_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 instr[5] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput24 read_data[15] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_204_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput35 start net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout110_I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3460_ _1149_ _1136_ _1152_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout208_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _2092_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3391_ _1045_ _1100_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2713__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5195__RN net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ _0292_ net206 clknet_leaf_88_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _0223_ net173 clknet_leaf_99_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_238_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4012_ _1530_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4769__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ _0076_ net282 clknet_leaf_31_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _0047_ net299 clknet_leaf_35_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_205_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4776_ _2142_ _0753_ _0714_ _2119_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_222_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3727_ _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3658_ _2169_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2609_ _2296_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4853__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3589_ _1161_ _1246_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5186__RN net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5328_ _0490_ net319 clknet_leaf_54_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5259_ _0421_ net236 clknet_leaf_72_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4457__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5209__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3004__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4209__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5359__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3939__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2843__I _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5110__RN net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_227_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4696__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4924__RN net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout190 net203 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2960_ net26 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout158_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5101__RN net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2891_ net79 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout325_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4630_ _1895_ _1965_ _1968_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4561_ _1923_ _1921_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2934__A1 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3512_ net25 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4492_ _2170_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3443_ _1127_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ _1021_ _1091_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5113_ _0275_ net205 clknet_leaf_88_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _0206_ net102 clknet_leaf_109_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_239_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5340__RN net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4611__A1 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _0030_ net148 clknet_leaf_17_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_194_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4759_ _1004_ _2046_ _2049_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3494__I _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2925__A1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5159__RN net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5031__CLK clknet_leaf_67_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4906__RN net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3102__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_50_clk_I clknet_4_13_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4899__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_223_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3169__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2916__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_65_clk_I clknet_4_12_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2519__I1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3090_ _0884_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3644__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3992_ _1529_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_18_clk_I clknet_4_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2943_ _0570_ _0773_ _0727_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2874_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4613_ _1927_ _1954_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5054__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4544_ _0603_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3580__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _1840_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3426_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout90_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3332__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3357_ _0991_ _1078_ _1082_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3288_ _1035_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _0189_ net105 clknet_leaf_118_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_227_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3489__I _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3399__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3571__A1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3952__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output71_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2568__I _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5077__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4023__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2590_ _2159_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3562__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ _1699_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4914__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2478__I _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3211_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4191_ _1633_ _1664_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3865__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3142_ _0921_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3073_ _0595_ _0606_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3617__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3975_ _1378_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4042__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2926_ Control_unit2.instr_stage2\[10\] _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_206_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2857_ _0696_ _0697_ net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2788_ Stack_pointer.SP\[1\] _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4527_ _1895_ _1891_ _1897_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4458_ _1742_ _1847_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2388__I _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3409_ _1058_ _1112_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4389_ _1780_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4281__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2595__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4937__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3544__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3682__I _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4272__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4024__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout140_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _1352_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout238_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0570_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3783__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3691_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2642_ _2323_ _2327_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5361_ _0523_ net139 clknet_leaf_21_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2573_ _2250_ _2095_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _1748_ _1739_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5292_ _0454_ net199 clknet_leaf_67_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ _1642_ _1700_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3838__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4174_ _1609_ _1655_ _1657_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_210_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3125_ _0591_ _0905_ _0908_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_228_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2936__I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_228_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3056_ _0824_ _2337_ _0856_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4263__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3958_ _1456_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2909_ net58 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3889_ _1446_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4254__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_203_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_226_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3677__I _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5115__CLK clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5265__CLK clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_4_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A2 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout188_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4930_ _0092_ net266 clknet_leaf_25_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout355_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ Stack_pointer.SP_next\[5\] net115 clknet_leaf_8_clk Stack_pointer.SP\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3056__I0 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3812_ _1376_ _1403_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4792_ _2067_ _0731_ _2073_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_221_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3743_ _1360_ _1356_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3674_ _1204_ _1302_ _1305_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2625_ _2226_ _2227_ _2243_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5344_ _0506_ net324 clknet_leaf_53_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4181__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2556_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5275_ _0437_ net236 clknet_leaf_68_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2487_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[2\].i3 _2110_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _1670_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2495__A1 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ _1201_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3108_ _0808_ _0894_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4088_ _1592_ _1586_ _1593_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4236__A2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3039_ _0798_ _2205_ _0842_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2798__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3995__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3497__I _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3047__I0 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3747__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__CLK clknet_leaf_116_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_112_clk clknet_4_0_0_clk clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2707__C1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5288__CLK clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout350 net351 net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2486__A1 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput14 instr[6] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput25 read_data[1] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_103_clk clknet_4_9_0_clk clknet_leaf_103_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_156_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2410_ _2092_ _2096_ _2100_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_196_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout103_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3390_ _0977_ _1098_ _1103_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_237_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3870__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _0222_ net180 clknet_leaf_103_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4011_ _1465_ _1538_ _1543_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3977__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4913_ _0075_ net282 clknet_leaf_30_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4206__I _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3110__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4844_ _0046_ net297 clknet_leaf_37_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _2058_ _0732_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3726_ _0614_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5184__D _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3657_ _1285_ _1289_ _1292_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2608_ _2279_ _2284_ _2295_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_162_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3588_ _1153_ _1245_ _1247_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2539_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5327_ _0489_ net317 clknet_leaf_53_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_5607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _0420_ net200 clknet_leaf_68_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input33_I read_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4209_ _1648_ _1678_ _1680_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5189_ _0351_ net161 clknet_leaf_98_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4209__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4116__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3955__I _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3196__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3690__I _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2459__A1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[1\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout180 net184 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout191 net195 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5303__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3959__A1 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2890_ Control_unit2.instr_stage2\[5\] _0713_ _0727_ _2273_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_203_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4560_ net25 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4384__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout318_I net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ _1123_ _1189_ _1194_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4491_ _1864_ _1867_ _1870_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3442_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4687__A2 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3373_ _1014_ _1090_ _1092_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _0274_ net168 clknet_leaf_92_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _0205_ net102 clknet_leaf_108_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_230_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_226_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_240_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4827_ _0029_ net147 clknet_leaf_19_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[4\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4820__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ _0815_ _2047_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ _0569_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4689_ _2004_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4970__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_12_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2689__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5326__CLK clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3015__I _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4602__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5095__RN net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4842__RN net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3685__I _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2764__I _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout170_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2852__A1 Control_unit2.instr_stage2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout268_I net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3991_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4843__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2942_ _2089_ _0712_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_200_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3595__I _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2873_ _0667_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4357__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_198_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4612_ _1873_ _1952_ _1957_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4993__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4543_ _1907_ _1903_ _1909_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4474_ _1838_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3425_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3332__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3356_ _0992_ _1079_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_213_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5010__RN net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout83_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3287_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _0188_ net105 clknet_leaf_118_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3096__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92_clk clknet_4_8_0_clk clknet_leaf_92_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_246_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5077__RN net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4824__RN net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4348__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3020__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output64_I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3087__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2584__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2834__A1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_83_clk clknet_4_10_0_clk clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5068__RN net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3562__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3210_ _2170_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4190_ _1629_ _1663_ _1667_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3141_ _2084_ _2135_ _2163_ _2185_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_6480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3072_ _0608_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_209_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3078__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_74_clk clknet_4_11_0_clk clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_236_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4578__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5059__RN net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3974_ _1476_ _1514_ _1519_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2925_ _2341_ _2352_ _0727_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4806__RN net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2856_ Control_unit1.instr_stage1\[6\] _0672_ _0684_ Stack_pointer.SP\[6\] _0697_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__CLK clknet_leaf_113_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2787_ _0620_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4750__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4526_ _1896_ _1893_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3553__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2669__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4457_ _1789_ _1846_ _1848_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3408_ _1005_ _1111_ _1114_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4388_ _1777_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3339_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3069__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _0171_ net108 clknet_leaf_107_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2816__A1 Stack_pointer.SP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_64_clk_I clknet_4_12_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_65_clk clknet_4_12_0_clk clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_79_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3241__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4741__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5222__RN net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_17_clk_I clknet_4_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4794__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2807__A1 Stack_pointer.SP\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_56_clk clknet_4_14_0_clk clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5044__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_233_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4034__I _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_0_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2710_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout133_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3783__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ _2321_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2641_ _2324_ _2326_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3873__I _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout300_I net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2572_ _2230_ _2260_ _2239_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5360_ _0522_ net323 clknet_leaf_53_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ net31 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5291_ _0453_ net236 clknet_leaf_72_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4242_ _1583_ _1698_ _1701_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3299__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ _1611_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3124_ _0832_ _0906_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3055_ _2338_ _0844_ _0858_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_215_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_47_clk clknet_4_15_0_clk clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_209_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_227_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_224_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3471__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2952__I _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3957_ _1498_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2908_ net58 _0742_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3888_ _1137_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2839_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4723__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5204__RN net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _1881_ _1877_ _1883_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_219_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5067__CLK clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4119__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3023__I _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_clk clknet_4_13_0_clk clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4904__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3693__I _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4714__A1 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4190__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_29_clk clknet_4_13_0_clk clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout250_I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4860_ Stack_pointer.SP_next\[4\] net116 clknet_leaf_8_clk Stack_pointer.SP\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA_fanout348_I net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3811_ _1325_ _1402_ _1405_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4791_ _0688_ _0668_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3056__I1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3742_ _1198_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3673_ _1303_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4705__A1 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2624_ _2265_ _2287_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_220_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _0505_ net323 clknet_leaf_53_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4181__A2 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2555_ _2236_ _2241_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_66_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5274_ _0436_ net200 clknet_leaf_69_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2486_ _2162_ _2146_ _2147_ _2178_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4225_ _1661_ _1684_ _1689_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_214_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4156_ _1592_ _1637_ _1645_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_229_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3107_ _2277_ _0893_ _0897_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4087_ _1503_ _1588_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_209_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3038_ _2192_ _0843_ _0848_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3444__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3995__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3047__I1 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4989_ _0151_ net315 clknet_leaf_56_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3747__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4402__I _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2707__B1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2707__C2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3018__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout340 net345 net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout351 net352 net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2486__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3435__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3738__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput15 instr[7] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput26 read_data[2] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2410__A2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5232__CLK clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5382__CLK clknet_leaf_28_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4010_ _1466_ _1539_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3674__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4912_ _0074_ net350 clknet_leaf_44_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_185_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4843_ _0045_ net287 clknet_leaf_32_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_209_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3729__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ net47 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2937__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3725_ _1344_ _1335_ _1346_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_clk clknet_4_5_0_clk clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3656_ _1191_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2607_ _2279_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3587_ _1156_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5326_ _0488_ net316 clknet_leaf_56_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2538_ _2225_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _0419_ net232 clknet_leaf_72_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2469_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4208_ _1597_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5188_ _0350_ net80 clknet_leaf_113_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_151_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input26_I read_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4139_ _1347_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4393__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4132__I _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_234_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2459__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout170 net171 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3656__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout181 net184 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_208_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout192 net195 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_208_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4307__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3211__I _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3959__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_231_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3510_ _1191_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout213_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4490_ _1779_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3441_ net28 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3881__I _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3372_ _1016_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2497__I _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ _0273_ net167 clknet_leaf_95_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ _0204_ net102 clknet_leaf_108_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3647__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5128__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4217__I _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3121__I _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5278__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2622__A2 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2960__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4826_ _0028_ net133 clknet_leaf_19_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[3\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4375__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _0998_ _2046_ _2048_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_198_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3708_ _1218_ _1320_ _1332_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4688_ _0933_ _1286_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3639_ _1260_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3886__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5309_ _0471_ net315 clknet_leaf_59_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_5416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4127__I _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4063__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3966__I _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_235_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4118__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3877__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3206__I _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2852__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout163_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2941_ _0712_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout330_I net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2872_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ _1925_ _1954_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ _1908_ _1905_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4473_ _1802_ _1852_ _1857_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3424_ _0879_ _0933_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3355_ _0987_ _1078_ _1081_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2540__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2540__B2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3286_ _1031_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5025_ _0187_ net186 clknet_leaf_106_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3052__S _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3096__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4596__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4809_ _0011_ net286 clknet_leaf_34_clk net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4348__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3859__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2531__B2 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output57_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3087__A2 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_233_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2598__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2598__B2 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4339__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2770__A1 Control_unit1.instr_stage1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3140_ _2205_ _2273_ _2251_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_6470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2775__I _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout280_I net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3071_ _0610_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4960__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3973_ _1518_ _1515_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_245_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2924_ _0751_ _0731_ _0757_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2855_ Control_unit2.instr_stage2\[6\] _0679_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5316__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2786_ Stack_pointer.SP\[1\] _0622_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4525_ net33 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4456_ _1738_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4990__RN net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3407_ _1006_ _1112_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _1802_ _1796_ _1803_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_219_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3269_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5008_ _0170_ net318 clknet_leaf_55_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2752__A1 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4140__I _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4981__RN net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4833__CLK clknet_4_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_5087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5339__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__I _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout126_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _2317_ _2305_ _2325_ _2307_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2571_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4310_ _1314_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_236_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5290_ _0452_ net194 clknet_leaf_69_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4241_ _1638_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_206_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4496__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4172_ _1639_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3123_ _0571_ _0905_ _0907_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4248__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3054_ _0818_ _0842_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_208_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3956_ _1495_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2907_ _0737_ _0738_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_220_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3887_ _1444_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2982__A1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2838_ _0616_ _0667_ _0675_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4856__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__A2 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2769_ Control_unit1.instr_stage1\[0\] _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2734__A1 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4508_ _1882_ _1879_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4439_ _1774_ _1832_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__B _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3304__I _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__RN net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4135__I _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_230_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_243_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5011__CLK clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3214__I _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5161__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2661__B1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__I _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3810_ _1326_ _1403_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout243_I net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4790_ _2189_ _0754_ _0733_ _2071_ _0709_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_162_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ _1294_ _1353_ _1359_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3884__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3672_ _1290_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2623_ _2299_ _2303_ _2309_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5198__RN net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_63_clk_I clknet_4_12_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2716__B2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5342_ _0504_ net323 clknet_leaf_53_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2554_ _2226_ _2227_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5273_ _0435_ net231 clknet_leaf_71_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2485_ _2083_ _2177_ _2099_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _1619_ _1685_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_78_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3141__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _1644_ _1640_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5370__RN net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3106_ _0805_ _0894_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4086_ _1296_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3037_ _0791_ _0842_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3060__S _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__RN net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_clk_I clknet_4_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _0150_ net311 clknet_leaf_59_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3939_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2955__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5189__RN net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2707__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2707__B2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5034__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout330 net332 net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout341 net345 net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3132__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout352 net353 net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__CLK clknet_leaf_87_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2486__A3 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4632__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput16 instr[8] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput27 read_data[3] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_204_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout193_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4623__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4911_ _0073_ net349 clknet_leaf_44_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_234_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4842_ _0044_ net285 clknet_leaf_33_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4773_ _1027_ _2052_ _2057_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_222_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2937__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4503__I _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5057__CLK clknet_leaf_103_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3724_ _1345_ _1337_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ _2287_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3586_ _1233_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4918__RN net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5325_ _0487_ net316 clknet_leaf_59_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_216_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2537_ _2226_ _2227_ _2223_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5256_ _0418_ net196 clknet_leaf_105_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2468_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[2\].i3 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_192_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3114__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _1672_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5187_ _0349_ net80 clknet_leaf_112_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2399_ _2080_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3665__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4138_ _1629_ _1622_ _1631_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input19_I read_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ _1486_ _1578_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_244_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__SETN net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3417__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4614__A1 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2928__A1 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3353__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout160 net166 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout171 net172 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout182 net184 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout193 net195 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3699__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3592__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3440_ _1125_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout206_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4917__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3344__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3371_ _1072_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5110_ _0272_ net157 clknet_leaf_95_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_152_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _0203_ net101 clknet_leaf_109_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3647__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5325__RN net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4072__A2 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _0027_ net133 clknet_leaf_19_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[2\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _0811_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3583__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3707_ _1331_ _1322_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4687_ _1913_ _1998_ _2003_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3638_ _1258_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3335__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3569_ _1196_ _1234_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3886__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5308_ _0470_ net199 clknet_leaf_62_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_5406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _0401_ net183 clknet_leaf_104_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5222__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4063__A2 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_223_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5372__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3574__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3877__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3222__I _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4054__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2940_ net50 _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_204_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3801__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2871_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout323_I net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _1871_ _1952_ _1956_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ net22 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3892__I _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4472_ _1760_ _1853_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3317__A1 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3423_ _0961_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3868__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3354_ _0988_ _1079_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2540__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3285_ _0930_ _1032_ _0759_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5245__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5024_ _0186_ net254 clknet_leaf_76_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2971__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4808_ _0010_ net285 clknet_leaf_34_clk net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3556__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _0973_ _2033_ _2037_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2531__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3042__I _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2881__I _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2598__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3795__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_197_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3547__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5118__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2830__B Control_unit1.instr_stage1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2770__A2 Control_unit1.instr_stage1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5268__CLK clknet_leaf_118_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3070_ _0864_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4275__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout273_I net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4027__A2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3887__I _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3972_ _1215_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2923_ _0752_ _0668_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_206_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2854_ _0694_ _0695_ net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3538__A1 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2785_ _0639_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4511__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4524_ _2335_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2761__A2 Arithmetic_Logic_Unit.ALU_001.p_Z vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ _1840_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3406_ _0999_ _1111_ _1113_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4386_ _1760_ _1797_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3337_ _1031_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3268_ _0590_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4266__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ _0169_ net318 clknet_leaf_55_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3199_ Control_unit2.instr_stage2\[10\] _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3797__I _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4833__D _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3529__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4421__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2752__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2876__I _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4257__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3768__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4331__I _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4193__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5090__CLK clknet_leaf_110_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2570_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout119_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _1699_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_218_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4496__A2 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4171_ _1636_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3122_ _0828_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4248__A2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3053_ _0857_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4506__I _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3955_ _1364_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4420__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2906_ _0737_ _0720_ _0711_ _0741_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3886_ _1453_ _1445_ _1454_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2837_ _0671_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3058__S _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2768_ Control_unit1.instr_stage1\[1\] _2115_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4507_ net29 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2699_ _2331_ _2380_ _2360_ _2381_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_191_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _1770_ _1831_ _1835_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4369_ _1789_ _1790_ _1792_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3320__I _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_208_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_115_clk clknet_4_0_0_clk clknet_leaf_115_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_210_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4151__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3990__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4950__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4478__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2489__A1 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5306__CLK clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2661__B2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_106_clk clknet_4_2_0_clk clknet_leaf_106_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_242_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3740_ _1358_ _1356_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout236_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3671_ _1137_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2622_ _2304_ _2308_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2716__A2 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2553_ _2223_ _2240_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5341_ _0503_ net321 clknet_leaf_51_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2484_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[2\].i3 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5272_ _0434_ net187 clknet_leaf_66_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4469__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4223_ _1617_ _1684_ _1688_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_229_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3141__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4154_ _1198_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3105_ _2256_ _0893_ _0896_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_233_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4085_ _1590_ _1586_ _1591_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3036_ _2177_ _0843_ _0847_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4641__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4987_ _0149_ net311 clknet_leaf_59_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_212_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4823__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3938_ _1186_ _1414_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_240_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3869_ _1348_ _1436_ _1441_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4973__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2707__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3380__A2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5329__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout320 net327 net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3315__I _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout331 net332 net331 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout342 net344 net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_232_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout353 net354 net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_232_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4146__I _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_243_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__RN net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 instr[9] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput28 read_data[4] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2410__A4 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3123__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout186_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4056__I _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ _0072_ net348 clknet_leaf_43_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout353_I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4841_ _0043_ net284 clknet_leaf_33_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4387__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4772_ _0837_ _2053_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4996__CLK clknet_4_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3723_ _1179_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3654_ _1287_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2605_ _2225_ _2241_ _2266_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3585_ _1231_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5324_ _0486_ net305 clknet_leaf_58_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__RN net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2536_ _2175_ _2196_ _2200_ _2218_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout99_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _0417_ net183 clknet_leaf_105_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2467_ _2132_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4206_ _1670_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2398_ Arithmetic_Logic_Unit.ALU_000.ALU_func\[0\] Arithmetic_Logic_Unit.ALU_000.ALU_func\[1\]
+ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_229_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5186_ _0348_ net80 clknet_leaf_112_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ _1630_ _1624_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_244_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _1480_ _1577_ _1579_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_225_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A2 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3019_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2625__A1 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4854__RN net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5001__CLK clknet_leaf_57_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2928__A2 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout150 net151 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout161 net165 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout172 net178 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4869__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2884__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout183 net184 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout194 net195 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_232_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5098__RN net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_clk_I clknet_4_12_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4845__RN net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__I _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4369__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5270__RN net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_221_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout101_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3370_ _1070_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5040_ _0202_ net255 clknet_leaf_76_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_clkbuf_leaf_15_clk_I clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2607__A1 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5089__RN net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5024__CLK clknet_leaf_76_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__RN net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4514__I _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4824_ _0026_ net133 clknet_leaf_19_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[1\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5174__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _2034_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3706_ _1165_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__RN net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4686_ _1914_ _1999_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2969__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3637_ _1218_ _1272_ _1277_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3335__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4532__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5013__RN net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3568_ _1123_ _1232_ _1235_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _0469_ net237 clknet_leaf_67_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2519_ _2203_ _2209_ _2210_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3499_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5238_ _0400_ net181 clknet_leaf_104_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input31_I read_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2846__A1 Control_unit2.instr_stage2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5169_ _0331_ net89 clknet_leaf_115_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_95_clk clknet_4_8_0_clk clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4827__RN net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4771__A1 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_86_clk clknet_4_10_0_clk clknet_leaf_86_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5047__CLK clknet_leaf_102_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5197__CLK clknet_leaf_83_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2870_ _2088_ _2090_ net35 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4762__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4540_ _0590_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout316_I net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10_clk clknet_4_5_0_clk clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4471_ _1758_ _1852_ _1856_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3317__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3422_ _1028_ _1117_ _1122_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3353_ _1047_ _1078_ _1080_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3284_ Control_unit2.instr_stage2\[9\] _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _0185_ net254 clknet_leaf_55_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3413__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_clk clknet_4_11_0_clk clknet_leaf_77_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_239_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _0009_ net285 clknet_leaf_34_clk net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_222_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2999_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4753__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3556__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ _0785_ _2035_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5234__RN net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4669_ _1980_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3323__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_68_clk clknet_4_9_0_clk clknet_leaf_68_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_245_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4907__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4154__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_198_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3795__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3993__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__RN net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3233__I _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_59_clk clknet_4_14_0_clk clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_236_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3235__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3971_ _1473_ _1514_ _1517_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2922_ _2335_ _0754_ _0733_ _0755_ _0710_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_210_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2853_ Control_unit1.instr_stage1\[5\] _0683_ _0685_ Stack_pointer.SP\[5\] _0695_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5216__RN net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2784_ _0627_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _1890_ _1891_ _1894_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5212__CLK clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4454_ _1838_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3405_ _1001_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4385_ _1378_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3336_ _0747_ _0752_ _0963_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5362__CLK clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4239__I _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3267_ _1014_ _1015_ _1018_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _0168_ net315 clknet_leaf_55_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3474__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3198_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3226__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3777__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2423__S _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4702__I _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__RN net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output62_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3988__I _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3217__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4193__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3228__I _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4170_ _1606_ _1649_ _1654_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3121_ _0887_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3052_ _0816_ _2318_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3208__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3954_ _1453_ _1496_ _1506_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2905_ Control_unit2.instr_stage2\[7\] _0713_ _0707_ _2272_ _0740_ _0741_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3885_ _1362_ _1447_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4708__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2836_ _2084_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2767_ Control_unit1.instr_decoder1.A\[0\] Control_unit1.instr_stage1\[2\] _0623_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4506_ _2255_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2698_ _2359_ _2358_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2977__I _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _1771_ _1832_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4368_ _1738_ _1791_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3319_ _1005_ _1054_ _1057_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4299_ _1728_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5108__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_230_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2422__A2 Control_unit1.instr_stage1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4432__I _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4175__A2 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3438__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3989__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3610__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout131_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout229_I net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3670_ _1288_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2621_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i2 _2305_ _2306_ _2307_ _2308_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4166__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5340_ _0502_ net274 clknet_leaf_61_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2552_ _2236_ _2225_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3913__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5271_ _0433_ net196 clknet_leaf_66_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2483_ _2128_ _2172_ _2175_ _2151_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4222_ _1659_ _1685_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4153_ _1590_ _1637_ _1643_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_228_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3104_ _0802_ _0894_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3429__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4084_ _1501_ _1588_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_244_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3035_ _0788_ _0844_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_209_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4986_ _0148_ net307 clknet_leaf_59_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3937_ _1491_ _1481_ _1493_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3601__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3868_ _1349_ _1437_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2819_ _0618_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3799_ _1365_ _1396_ _1398_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout310 net313 net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout321 net326 net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3668__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout332 net339 net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout343 net344 net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout354 net355 net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5080__CLK clknet_leaf_101_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4396__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4162__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 read_data[0] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 read_data[5] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3506__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4337__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout179_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout346_I net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _0042_ net287 clknet_leaf_32_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4771_ _1023_ _2052_ _2056_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3722_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3653_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2604_ _2246_ _2289_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_122_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3584_ _1149_ _1239_ _1244_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5323_ _0485_ net304 clknet_leaf_57_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2535_ _2120_ _2127_ _2214_ _2215_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_170_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5254_ _0416_ net181 clknet_leaf_104_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2466_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4205_ _1594_ _1671_ _1677_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5185_ _0347_ net89 clknet_leaf_113_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2397_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[0\].i3 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ _1179_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ _1482_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3018_ net23 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2625__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2990__I _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4940__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _0131_ net331 clknet_leaf_40_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_145_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4550__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3326__I _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout140 net141 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout151 net152 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout162 net165 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout173 net174 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_219_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout184 net190 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_235_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout195 net202 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2864__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4157__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3813__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4813__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_207_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4963__CLK clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _0025_ net133 clknet_leaf_3_clk Arithmetic_Logic_Unit.ALU_001.Y_CY\[0\].i3
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4754_ _2032_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3705_ _1329_ _1320_ _1330_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _1910_ _1998_ _2002_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2791__A1 Stack_pointer.SP\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3636_ _1166_ _1273_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3567_ _1191_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5306_ _0468_ net273 clknet_leaf_62_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2518_ _2159_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_192_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3498_ net24 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2985__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5237_ _0399_ net182 clknet_leaf_104_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2449_ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3099__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _0330_ net219 clknet_leaf_86_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2846__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input24_I read_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4119_ _1328_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4048__A1 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5099_ _0261_ net212 clknet_leaf_91_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_217_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4599__A2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3271__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4771__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2534__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4986__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4615__I _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4762__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2773__A1 Stack_pointer.SP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout211_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4350__I _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout309_I net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ _1800_ _1853_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3421_ _1029_ _1118_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2525__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3352_ _0983_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3283_ _0932_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5022_ _0184_ net250 clknet_leaf_75_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5141__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4450__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _0008_ net121 clknet_leaf_13_clk net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4202__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2998_ net19 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ _0961_ _2033_ _2036_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4260__I _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4668_ _1978_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4993__RN net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3619_ _1260_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4599_ _1910_ _1944_ _1948_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_61_clk_I clknet_4_12_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_76_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__A1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_14_clk_I clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4984__RN net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_29_clk_I clknet_4_13_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5014__CLK clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3180__A1 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5164__CLK clknet_leaf_90_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4345__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout161_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3970_ _1474_ _1515_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout259_I net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2921_ net59 _0743_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_182_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2852_ Control_unit2.instr_stage2\[5\] _0681_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2783_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4080__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _1892_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4453_ _1735_ _1839_ _1845_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_236_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3404_ _1099_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4384_ _1758_ _1796_ _1801_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_217_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3171__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3335_ _1028_ _1062_ _1067_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3266_ _1016_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5005_ _0167_ net315 clknet_leaf_56_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3197_ _2143_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3474__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4671__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4726__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4966__RN net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3162__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5187__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output55_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5143__RN net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4414__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3509__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3244__I _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3120_ _0885_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3051_ _0850_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4653__A1 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5134__RN net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4075__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4405__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3953_ _1505_ _1499_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2904_ _0732_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3884_ _1299_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ _0678_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2766_ _0620_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3392__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4505_ _1789_ _1877_ _1880_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2697_ _2337_ _2259_ _2357_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4436_ _1767_ _1831_ _1834_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3144__A1 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ _1780_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5373__RN net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3318_ _1006_ _1055_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4298_ net28 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3249_ _2335_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5125__RN net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2958__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4939__RN net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3135__A1 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5116__RN net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2661__A3 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5202__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3239__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2620_ _2149_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout124_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2551_ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_182_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5270_ _0432_ net185 clknet_leaf_106_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2482_ _2174_ _2151_ _2154_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__3126__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_233_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4221_ _1614_ _1684_ _1687_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5355__RN net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4152_ _1642_ _1640_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3141__A4 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3103_ _0795_ _0893_ _0895_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2519__S _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4083_ _1293_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3702__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3034_ _2148_ _0843_ _0846_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_243_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4985_ _0147_ net307 clknet_leaf_59_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3936_ _1492_ _1483_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3601__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _1344_ _1436_ _1440_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2818_ _0638_ _0640_ _0664_ _0666_ Stack_pointer.SP_next\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_3798_ _1303_ _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2988__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2749_ _0561_ _0562_ _0581_ _0597_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout300 net301 net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4419_ _1748_ _1820_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout311 net313 net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout322 net326 net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout333 net338 net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout344 net345 net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout355 net34 net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_232_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5225__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4443__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_230_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 read_data[10] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3356__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_237_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3108__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4608__A1 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4353__I _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout241_I net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout339_I net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _0834_ _2053_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ _0603_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3652_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3347__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2603_ _2290_ _2266_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4892__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3583_ _1151_ _1240_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3898__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2534_ _2216_ _2219_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5322_ _0484_ net304 clknet_leaf_58_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2465_ _2140_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _0415_ net187 clknet_leaf_65_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5248__CLK clknet_leaf_77_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4204_ _1646_ _1673_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5184_ _0346_ net218 clknet_leaf_87_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2396_ _2091_ net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4528__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4135_ _1343_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4066_ _1559_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3017_ _0591_ _0826_ _0833_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_168_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3822__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4968_ _0130_ net293 clknet_leaf_38_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_196_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3919_ _1379_ _1469_ _1479_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4899_ _0061_ net285 clknet_leaf_33_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3607__I _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout130 net132 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2667__B _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout141 net142 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout152 net153 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3510__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout163 net165 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout174 net177 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_232_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout185 net189 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout196 net201 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_235_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_228_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3577__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3517__I _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__A2 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3501__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout191_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout289_I net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4057__A2 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4083__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4822_ _0024_ net347 clknet_leaf_44_clk net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_221_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3568__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4753_ _0994_ _2040_ _2045_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ _1216_ _1322_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4684_ _1911_ _1999_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ _1163_ _1272_ _1276_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5305_ _0467_ net304 clknet_leaf_62_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3740__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2517_ _2161_ _2185_ _2205_ _2207_ _2208_ _2163_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_192_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3497_ _1027_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2448_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5236_ _0398_ net100 clknet_leaf_111_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _0329_ net220 clknet_leaf_85_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4118_ _1614_ _1610_ _1616_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_244_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5098_ _0260_ net232 clknet_leaf_70_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4048__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input17_I instr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4049_ _1460_ _1566_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_244_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4721__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2534__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3731__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4039__A2 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4211__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5093__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _1024_ _1117_ _1121_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout204_I net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2525__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3351_ _1072_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3282_ _1028_ _1015_ _1030_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4278__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I instr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _0183_ net249 clknet_leaf_74_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4078__I _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3710__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2461__A1 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4805_ _0007_ net121 clknet_leaf_13_clk net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_206_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2997_ _2336_ _0810_ _0817_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_222_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4202__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4541__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _0780_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3157__I _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _1887_ _1986_ _1991_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3618_ _1258_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4598_ _1911_ _1945_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3549_ _1192_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5219_ _0381_ net81 clknet_leaf_112_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4441__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_205_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3067__I _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4953__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3704__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5309__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4680__A2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4626__I _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2691__B2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2920_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout154_I net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2851_ _0692_ _0693_ net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_223_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout321_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2782_ _0626_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4521_ _1868_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ _1787_ _1841_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A2 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3403_ _1097_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_236_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4383_ _1800_ _1797_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3334_ _1029_ _1063_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3265_ _0970_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _0166_ net307 clknet_leaf_56_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3196_ _0615_ _0955_ _0960_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4536__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3440__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4826__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4976__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4719_ _0823_ _2020_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_202_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3162__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output48_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2673__A1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3350__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4414__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2425__A1 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_118_clk clknet_4_1_0_clk clknet_leaf_118_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5131__CLK clknet_leaf_89_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3525__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2900__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5281__CLK clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3050_ _0855_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4849__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4653__A2 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout271_I net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4356__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2664__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4893__RN net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_109_clk clknet_4_0_0_clk clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_60_clk_I clknet_4_12_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3952_ _1201_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4999__CLK clknet_leaf_63_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2903_ net57 _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3883_ _1451_ _1445_ _1452_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2834_ _0633_ _0677_ _0680_ net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2719__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_75_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3916__A1 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2765_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _1878_ _1879_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5070__RN net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2696_ _2299_ _2303_ _2378_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_201_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4435_ _1768_ _1832_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3144__A2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4366_ _1777_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3317_ _0999_ _1054_ _1056_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4297_ _1726_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_clk_I clknet_4_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3248_ _0999_ _1000_ _1003_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2495__B _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4644__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2655__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3179_ _0812_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2655__B2 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_215_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_28_clk_I clknet_4_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5004__CLK clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5061__RN net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_237_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3135__A2 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4875__RN net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__I _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3374__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout117_I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2550_ _2237_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3255__I _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2481_ _2092_ _2173_ _2100_ _2104_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3126__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4220_ _1615_ _1685_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _1195_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2885__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3102_ _0798_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _1583_ _1586_ _1589_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4086__I _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3033_ _0785_ _0844_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2637__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5027__CLK clknet_leaf_118_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__RN net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _0146_ net272 clknet_leaf_63_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5177__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3935_ _1183_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__RN net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3866_ _1345_ _1437_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2817_ Control_unit1.instr_stage1\[10\] _0637_ _0639_ _0664_ _0665_ _0666_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_165_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3797_ _1390_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4562__A1 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2748_ _0576_ _0597_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_219_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2679_ _2358_ _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4418_ _1744_ _1819_ _1823_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout301 net302 net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout312 net313 net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_207_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout323 net324 net323 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout334 net338 net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4349_ _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout345 net350 net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4871__D Control_unit1.instr_stage1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4608__A2 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2419__I Control_unit1.instr_decoder1.A\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2619__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3292__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3720_ _1340_ _1335_ _1342_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout234_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_40_clk clknet_4_15_0_clk clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_187_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3651_ _1229_ _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3347__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2602_ _2230_ _2235_ _2239_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_220_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3582_ _1145_ _1239_ _1243_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5321_ _0483_ net304 clknet_leaf_58_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2533_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5252_ _0414_ net106 clknet_leaf_108_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2464_ _2155_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_170_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4203_ _1592_ _1671_ _1676_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_218_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5183_ _0345_ net226 clknet_leaf_84_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3713__I _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2395_ _2088_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4134_ _1626_ _1622_ _1628_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4065_ _1557_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3016_ _0832_ _0829_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_225_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__RN net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4544__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3035__A1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4967_ _0129_ net293 clknet_leaf_29_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4783__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3918_ _1478_ _1471_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5264__RN net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_clk clknet_4_6_0_clk clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4898_ _0060_ net289 clknet_leaf_33_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2999__I _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3849_ _1315_ _1424_ _1429_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4866__D Control_unit1.instr_stage1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2849__A1 Control_unit2.instr_stage2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout120 net121 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xclkbuf_leaf_98_clk clknet_4_8_0_clk clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_232_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout142 net152 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout153 net154 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout164 net165 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout175 net177 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout186 net189 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5342__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout197 net201 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_210_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4454__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_22_clk clknet_4_2_0_clk clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3329__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__RN net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2552__A3 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_89_clk clknet_4_10_0_clk clknet_leaf_89_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_215_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3501__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout184_I net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout351_I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _0023_ net347 clknet_leaf_44_clk net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4752_ _0807_ _2041_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_226_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_13_clk clknet_4_4_0_clk clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_222_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3703_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ _1907_ _1998_ _2001_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4517__A1 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3634_ _1216_ _1273_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5215__CLK clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3565_ _1230_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _0466_ net188 clknet_leaf_65_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2516_ _2165_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3740__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout97_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3496_ _1178_ _1169_ _1181_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5365__CLK clknet_leaf_28_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5235_ _0397_ net94 clknet_leaf_111_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2447_ _2129_ _2139_ _2141_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3443__I _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5166_ _0328_ net226 clknet_leaf_84_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4117_ _1615_ _1612_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5097_ _0259_ net193 clknet_leaf_101_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ _1507_ _1565_ _1567_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3256__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_240_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4756__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3618__I _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3731__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3495__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4882__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4184__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__CLK clknet_leaf_104_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3350_ _1070_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2930__B1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4359__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3281_ _1029_ _1017_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3263__I _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _0182_ net238 clknet_leaf_73_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_239_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_2_clk clknet_4_6_0_clk clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3486__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3789__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2461__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4804_ _0006_ net119 clknet_leaf_5_clk net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4738__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ _0816_ _0813_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_222_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3410__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4666_ _1888_ _1987_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3961__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3617_ _1134_ _1259_ _1265_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4597_ _1907_ _1944_ _1947_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3548_ _1188_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4269__I _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3479_ _1060_ _1154_ _1167_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5218_ _0380_ net81 clknet_leaf_112_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5149_ _0311_ net217 clknet_leaf_87_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3901__I _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4729__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3401__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2507__A3 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2691__A2 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2427__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5060__CLK clknet_leaf_103_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2850_ Control_unit1.instr_stage1\[4\] _0683_ _0685_ Stack_pointer.SP\[4\] _0693_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout147_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2781_ Stack_pointer.SP\[1\] _0621_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3258__I _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ net32 _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout314_I net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4451_ _1733_ _1839_ _1844_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3402_ _0995_ _1105_ _1110_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4382_ net19 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_236_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3333_ _1024_ _1062_ _1066_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3264_ _0827_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3459__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _0165_ net306 clknet_leaf_57_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3195_ _0838_ _0956_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3721__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2434__A2 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3631__A1 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4187__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2979_ _2256_ _0796_ _0803_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3168__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4718_ _1008_ _2019_ _2023_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4649_ _1980_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4874__D Control_unit1.instr_stage1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5083__CLK clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2425__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3622__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4178__A2 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3925__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3806__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_214_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2866__B Arithmetic_Logic_Unit.ALU_001.p_Z vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3541__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout264_I net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _1451_ _1496_ _1504_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2416__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3613__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2902_ net55 net56 _0723_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_147_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3882_ _1360_ _1447_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2833_ _2079_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4169__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3916__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2764_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _1868_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2695_ _2329_ _2377_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3716__I _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2620__I _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4434_ _1762_ _1831_ _1833_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_236_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4365_ _1364_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3316_ _1001_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4296_ _1735_ _1727_ _1736_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3247_ _1001_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3451__I _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3178_ _0937_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2655__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4943__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3604__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__D Control_unit1.instr_stage1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_198_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output60_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3361__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4096__A1 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4020__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3536__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2480_ _2107_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4816__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_229_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4150_ _1583_ _1637_ _1641_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3101_ _0887_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4367__I _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4081_ _1497_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4087__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4966__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3032_ _2097_ _0843_ _0845_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2637__A2 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3834__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4983_ _0145_ net271 clknet_leaf_61_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3934_ _1347_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3865_ _1340_ _1436_ _1439_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2816_ Stack_pointer.SP\[7\] _0657_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ _1388_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2747_ _0604_ net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4562__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3446__I _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2678_ _2349_ _2350_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4417_ _1745_ _1820_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout302 net303 net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout313 net314 net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout324 net326 net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4348_ _0883_ _1186_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout335 net336 net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout346 net348 net346 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4279_ _1284_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5121__CLK clknet_leaf_98_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5271__CLK clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2564__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4305__A2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4989__CLK clknet_leaf_56_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3091__I _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2619__A2 Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_74_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_89_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4792__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3650_ _0747_ _1032_ _0759_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_201_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout227_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_12_clk_I clknet_4_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2601_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_228_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3581_ _1147_ _1240_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2555__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ _0482_ net188 clknet_leaf_65_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2532_ _2220_ _2222_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_196_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5251_ _0413_ net95 clknet_leaf_117_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2463_ _2156_ _2128_ _2105_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_27_clk_I clknet_4_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4202_ _1644_ _1673_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _0344_ net223 clknet_leaf_82_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2394_ _2089_ Control_unit2.instr_stage2\[11\] _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_233_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4097__I _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4133_ _1627_ _1624_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4064_ _1520_ _1571_ _1576_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_209_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5144__CLK clknet_leaf_93_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3015_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_225_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4966_ _0128_ net291 clknet_leaf_29_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__CLK clknet_leaf_74_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3917_ _1165_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_240_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4783__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4897_ _0059_ net287 clknet_leaf_32_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2794__A1 Control_unit1.instr_stage1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4560__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3848_ _1316_ _1425_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3779_ _1345_ _1382_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3904__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout110 net111 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout121 net127 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2849__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout132 net135 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout143 net144 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout154 net355 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout165 net166 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout176 net177 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout187 net189 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout198 net200 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4882__D net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4735__I _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4471__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3026__A2 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3086__I _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2537__A1 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5017__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5167__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5191__RN net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout177_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__C2 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4820_ _0022_ net346 clknet_leaf_44_clk net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout344_I net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3017__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4751_ _0990_ _2040_ _2044_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3702_ _2353_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4682_ _1908_ _1999_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3633_ _1159_ _1272_ _1275_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2528__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3564_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2515_ _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5303_ _0465_ net187 clknet_leaf_65_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3495_ _1180_ _1172_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2446_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _0396_ net93 clknet_leaf_111_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_237_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5165_ _0327_ net217 clknet_leaf_87_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_190_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5182__RN net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4116_ _1160_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5096_ _0258_ net177 clknet_leaf_100_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_244_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4047_ _1456_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4756__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4949_ _0111_ net292 clknet_leaf_37_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_166_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2767__A1 Control_unit1.instr_decoder1.A\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4996__RN net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4508__A2 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4877__D Control_unit1.instr_stage1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3495__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__RN net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4465__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4987__RN net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3183__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2930__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3280_ _0837_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout294_I net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4683__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3486__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__RN net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2997__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _0005_ net120 clknet_leaf_5_clk net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_222_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2995_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2749__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4734_ _2031_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _1884_ _1986_ _1990_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5332__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3616_ _1202_ _1261_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4596_ _1908_ _1945_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3547_ _1218_ _1211_ _1219_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2921__A1 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3478_ _1166_ _1157_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2429_ _2102_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5217_ _0379_ net89 clknet_leaf_114_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4674__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5155__RN net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _0310_ net213 clknet_leaf_90_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input22_I read_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4902__RN net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4285__I _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5079_ _0241_ net191 clknet_leaf_102_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4729__A2 _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3629__I _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3165__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5394__RN net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4665__A1 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4195__I _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__CLK clknet_leaf_99_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3640__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5355__CLK clknet_leaf_60_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2780_ _0628_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout307_I net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4450_ _1785_ _1841_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3401_ _0996_ _1106_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4381_ _1755_ _1796_ _1799_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3274__I _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2903__A1 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5385__RN net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3332_ _1025_ _1063_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3263_ _0968_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _0164_ net307 clknet_leaf_58_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3194_ _0604_ _0955_ _0959_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2618__I _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4408__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2978_ _0802_ _0799_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3395__A1 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _1940_ _2020_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4648_ _1977_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4872__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4579_ _1887_ _1930_ _1935_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5376__RN net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5128__RN net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__CLK clknet_leaf_101_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4890__D net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3386__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4638__A1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3310__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2438__I _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3950_ _1503_ _1499_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout257_I net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3613__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2901_ net57 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_205_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3269__I _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _1296_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2832_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3377__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4895__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2763_ _0616_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_185_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2901__I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4502_ net28 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2694_ _2347_ _2358_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_172_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4433_ _1764_ _1832_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5358__RN net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4364_ _1735_ _1778_ _1788_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3315_ _1038_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3732__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4295_ _1646_ _1729_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3246_ _0970_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3301__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3177_ _0935_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4563__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3604__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3368__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3907__I _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5050__CLK clknet_leaf_71_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2879__B1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__D net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3540__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output53_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3089__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3359__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3817__I _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4020__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3531__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3100_ _0885_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4080_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3031_ _0780_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2637__A3 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3834__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4982_ _0144_ net271 clknet_leaf_64_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3598__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3933_ _1488_ _1481_ _1490_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3864_ _1341_ _1437_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2815_ Stack_pointer.SP\[7\] _0620_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3795_ _1300_ _1389_ _1395_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3727__I _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5073__CLK clknet_leaf_104_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2746_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2573__A2 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2677_ _2331_ _2359_ _2360_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4416_ _1741_ _1819_ _1822_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5396_ _0558_ net120 clknet_leaf_11_clk net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout303 net353 net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3522__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout314 net328 net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout325 net326 net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3462__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4347_ _1773_ _1763_ _1775_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout336 net337 net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout347 net348 net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4910__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4278_ _1632_ _1717_ _1722_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_246_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3229_ _0801_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3825__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2806__I _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5096__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2451__I _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout122_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ _2250_ _2258_ _2264_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3052__I0 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3580_ _1141_ _1239_ _1242_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2555__A2 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2531_ _2204_ _2152_ _2221_ _2099_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ _0412_ net95 clknet_leaf_117_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4933__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2462_ _2112_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4201_ _1590_ _1671_ _1675_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2393_ Control_unit2.instr_stage2\[12\] _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5181_ _0343_ net213 clknet_leaf_83_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4132_ _1175_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _1478_ _1572_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3014_ net22 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4480__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4965_ _0127_ net293 clknet_leaf_29_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4232__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3916_ _1476_ _1469_ _1477_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4896_ net8 net144 clknet_leaf_16_clk Control_unit1.instr_decoder1.A\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3847_ _1311_ _1424_ _1428_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3457__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3043__I0 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3778_ _1340_ _1381_ _1384_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2546__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2729_ _0585_ _0566_ _0587_ _2207_ _2208_ _2365_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_173_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4288__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout100 net103 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5379_ _0541_ net268 clknet_leaf_25_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout111 net154 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout122 net126 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout133 net135 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout144 net145 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout155 net156 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout166 net179 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_232_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout177 net178 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout188 net189 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_210_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout199 net200 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_235_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_231_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4956__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2537__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3830__I _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_7_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2473__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2473__B2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout337_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4750_ _0804_ _2041_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3701_ _1325_ _1320_ _1327_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4681_ _1902_ _1998_ _2000_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3632_ _1161_ _1273_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2528__A2 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3563_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5302_ _0464_ net261 clknet_leaf_65_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2514_ _2136_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3494_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5111__CLK clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ _0395_ net100 clknet_leaf_108_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_170_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2445_ Arithmetic_Logic_Unit.op _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5164_ _0326_ net208 clknet_leaf_90_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2700__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4115_ _1324_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _0257_ net173 clknet_leaf_101_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ _1559_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4829__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4453__A2 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4205__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4571__I _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4948_ _0110_ net281 clknet_leaf_30_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4979__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2767__A2 Control_unit1.instr_stage1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3187__I _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4879_ Control_unit1.instr_decoder1.A\[1\] net143 clknet_leaf_16_clk Control_unit2.instr_decoder2.A\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_73_clk_I clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3192__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_88_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_11_clk_I clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_26_clk_I clknet_4_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3707__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__CLK clknet_leaf_85_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2930__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__CLK clknet_leaf_118_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4683__A2 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout287_I net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2694__A1 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4435__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4802_ _0004_ net119 clknet_leaf_5_clk net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2994_ net33 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4733_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _1885_ _1987_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3615_ _1132_ _1259_ _1264_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4595_ _1902_ _1944_ _1946_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3735__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3546_ _1166_ _1212_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3477_ _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4123__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5216_ _0378_ net223 clknet_leaf_83_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2428_ _2121_ _2122_ _2117_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4566__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5147_ _0309_ net208 clknet_leaf_89_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3470__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2685__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5078_ _0240_ net182 clknet_leaf_102_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input15_I instr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4426__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4029_ _1488_ _1550_ _1554_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5007__CLK clknet_leaf_55_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5091__RN net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3400_ _0991_ _1105_ _1109_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout202_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4380_ _1756_ _1797_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3331_ _1020_ _1062_ _1065_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3262_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I instr[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _0163_ net306 clknet_leaf_57_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3290__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3193_ _0835_ _0956_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4408__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3092__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3919__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2977_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4716_ _1004_ _2019_ _2022_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_206_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4647_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3465__I _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3147__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4578_ _1888_ _1931_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3529_ _1143_ _1206_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_15_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2745__S _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3083__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2544__I _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4583__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5064__RN net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2897__A1 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4638__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__RN net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5322__CLK clknet_leaf_58_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2454__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[1\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2900_ _0730_ _0731_ _0711_ _0736_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_225_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout152_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3880_ _1449_ _1445_ _1450_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_70_clk clknet_4_9_0_clk clknet_leaf_70_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_182_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2831_ _0616_ _2086_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3377__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5055__RN net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2762_ Control_unit2.instr_decoder2.A\[2\] _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2585__B1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4501_ _1866_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4802__RN net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2403__B Arithmetic_Logic_Unit.ALU_000.ALU_func\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2693_ _2375_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3129__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4326__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4432_ _1813_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4363_ _1787_ _1781_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3314_ _1035_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4294_ _1299_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3245_ _0811_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3176_ _2297_ _0943_ _0948_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_230_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2812__A1 Stack_pointer.SP\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5294__RN net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_61_clk clknet_4_12_0_clk clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_223_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4565__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2879__A1 Control_unit2.instr_stage2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3923__I _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2539__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5345__CLK clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output46_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4754__I _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2803__A1 Stack_pointer.SP\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5285__RN net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_52_clk clknet_4_14_0_clk clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_207_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput70 net70 write_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2449__I _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3030_ _0841_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3295__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4981_ _0143_ net271 clknet_leaf_61_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_224_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3598__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3932_ _1489_ _1483_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_43_clk clknet_4_15_0_clk clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_205_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3863_ _1334_ _1436_ _1438_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2912__I Control_unit2.instr_stage2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2814_ _0638_ _0640_ _0661_ _0663_ Stack_pointer.SP_next\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5218__CLK clknet_leaf_112_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3794_ _1362_ _1391_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _0599_ _0602_ _2249_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2676_ _2342_ _2347_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_219_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5368__CLK clknet_leaf_61_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4415_ _1742_ _1820_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5395_ _0557_ net122 clknet_leaf_11_clk net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout304 net308 net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5200__RN net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4346_ _1774_ _1765_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout315 net320 net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_236_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout326 net327 net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout337 net338 net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout348 net349 net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4277_ _1633_ _1718_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3228_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3159_ _0781_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A1 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_34_clk clknet_4_7_0_clk clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3139__B _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3653__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4710__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3277__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4885__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4484__I _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5258__RN net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_25_clk clknet_4_3_0_clk clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3828__I _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2732__I _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4529__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_224_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3052__I1 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_3_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout115_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2530_ _2130_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[4\].i3 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2888__B _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__I _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2461_ _2151_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_177_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ _1642_ _1673_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ _0342_ net211 clknet_leaf_91_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2392_ _2079_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4131_ _1339_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _1476_ _1571_ _1575_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3013_ _0571_ _0826_ _0830_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4768__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4964_ _0126_ net267 clknet_leaf_27_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_16_clk clknet_4_7_0_clk clknet_leaf_16_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5040__CLK clknet_leaf_76_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _1376_ _1471_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4895_ net7 net143 clknet_leaf_15_clk Control_unit1.instr_decoder1.A\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_205_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3846_ _1312_ _1425_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5190__CLK clknet_leaf_96_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3043__I1 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3777_ _1341_ _1382_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3743__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__I _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2659_ _2343_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3473__I _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5378_ _0540_ net268 clknet_leaf_26_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout101 net103 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout112 net113 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_216_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout123 net126 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout134 net135 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4329_ _1661_ _1751_ _1761_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout145 net151 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout156 net160 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout167 net168 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout178 net179 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3259__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout189 net190 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2482__A2 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4759__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3648__I _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3982__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2501__B _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3383__I _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__CLK clknet_leaf_100_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2473__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3422__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _1326_ _1322_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_187_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout232_I net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4680_ _1904_ _1999_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4900__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _1153_ _1272_ _1274_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_200_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3562_ _1226_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3725__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5301_ _0463_ net186 clknet_leaf_65_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2513_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4389__I _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3493_ net23 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5232_ _0394_ net225 clknet_leaf_84_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2444_ _2133_ _2106_ _2135_ _2137_ _2138_ _2118_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
Xclkbuf_leaf_5_clk clknet_4_4_0_clk clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5163_ _0325_ net209 clknet_leaf_89_clk net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4114_ _1609_ _1610_ _1613_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ _0256_ net182 clknet_leaf_103_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ _1557_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_212_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _0109_ net281 clknet_leaf_31_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3468__I _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3964__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4878_ Control_unit1.instr_decoder1.A\[0\] net143 clknet_leaf_15_clk Arithmetic_Logic_Unit.op
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4299__I _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4141__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3931__I _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5086__CLK clknet_leaf_78_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4380__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4002__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3841__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout182_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ _0003_ net119 clknet_leaf_12_clk net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4199__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2993_ _2322_ _0810_ _0814_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_210_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3288__I _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _2031_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4663_ _1881_ _1986_ _1989_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3614_ _1199_ _1261_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4594_ _1904_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3545_ _0821_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_200_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4371__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3476_ net20 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _0377_ net227 clknet_leaf_84_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2427_ net1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3751__I _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_213_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5146_ _0308_ net206 clknet_leaf_88_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5077_ _0239_ net163 clknet_leaf_99_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4946__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4028_ _1489_ _1551_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3634__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3198__I _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_4_11_0_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3937__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3926__I _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2676__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3625__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4492__I _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3928__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2600__A2 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__CLK clknet_leaf_117_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4819__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3330_ _1021_ _1063_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3261_ _0570_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _0162_ net273 clknet_leaf_63_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4969__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3192_ _0591_ _0955_ _0958_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3616__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_72_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2915__I _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3092__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_87_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3919__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2976_ net29 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4715_ _0815_ _2020_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2650__I _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4646_ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_10_clk_I clknet_4_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4577_ _1884_ _1930_ _1934_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3528_ _1204_ _1205_ _1207_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_25_clk_I clknet_4_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3481__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3459_ _1151_ _1139_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5129_ _0291_ net206 clknet_leaf_87_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5124__CLK clknet_leaf_116_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3083__A2 Control_unit2.instr_decoder2.A\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2560__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[6\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4335__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4487__I _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4099__A1 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2821__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2830_ _0672_ _0676_ Control_unit1.instr_stage1\[0\] _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout145_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2761_ _2140_ Arithmetic_Logic_Unit.ALU_001.p_Z _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3566__I _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2585__A1 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2585__B2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout312_I net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ _1875_ _1867_ _1876_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2692_ _2370_ _2374_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4431_ _1811_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4362_ net27 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3313_ _0995_ _1048_ _1053_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4293_ _1733_ _1727_ _1734_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3244_ _0968_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__CLK clknet_leaf_89_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3175_ _0808_ _0944_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5297__CLK clknet_leaf_118_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4565__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3476__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2959_ _2171_ _0779_ _0787_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_202_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4629_ _1896_ _1966_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4253__A1 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2803__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4005__A1 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput60 net60 write_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_218_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput71 net71 write_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout262_I net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4980_ _0142_ net262 clknet_leaf_24_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_184_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3931_ _1179_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _1336_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2813_ Control_unit1.instr_stage1\[9\] _0637_ _0639_ _0661_ _0662_ _0663_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4547__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3793_ _1297_ _1389_ _1394_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2744_ _0585_ _0587_ _0600_ _0601_ _2208_ _0566_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_185_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2675_ _2345_ _2346_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_201_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _1789_ _1819_ _1821_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5394_ _0556_ net124 clknet_leaf_14_clk net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout305 net308 net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4345_ net24 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_236_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout316 net320 net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2730__A1 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout327 net328 net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout338 net339 net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout349 net350 net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4276_ _1629_ _1717_ _1721_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_173_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3227_ _2255_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3286__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3158_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3089_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A2 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2797__A1 Stack_pointer.SP\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[5\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2549__B2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5312__CLK clknet_leaf_53_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3934__I _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4950__RN net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4765__I _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3277__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2788__A1 Stack_pointer.SP\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3201__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2460_ _2134_ _2096_ _2153_ _2150_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2391_ _2080_ Control_unit2.instr_decoder2.A\[1\] _2084_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__RN net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4130_ _1621_ _1622_ _1625_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4061_ _1518_ _1572_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3012_ _0828_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4768__A2 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _0125_ net267 clknet_leaf_27_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_224_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2779__A1 Stack_pointer.SP\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3914_ _1328_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4894_ net6 net146 clknet_leaf_15_clk Control_unit1.instr_decoder1.A\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_162_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5335__CLK clknet_leaf_64_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3845_ _1307_ _1424_ _1427_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3776_ _1334_ _1381_ _1383_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2727_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[14\].i3 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2658_ _2342_ _2331_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2589_ _2277_ net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5377_ _0539_ net268 clknet_leaf_26_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5185__RN net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout102 net103 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout113 net114 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_236_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2703__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout124 net126 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout135 net142 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4328_ _1760_ _1753_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout146 net147 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout157 net159 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout168 net172 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout179 net204 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4259_ _1697_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4456__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2482__A3 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3195__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4852__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4695__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5176__RN net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4923__RN net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4495__I _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5208__CLK clknet_leaf_97_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5358__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2743__I _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3422__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3630_ _1156_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout225_I net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3186__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3561_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _0462_ net104 clknet_leaf_119_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_183_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2512_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[4\].i3 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3492_ _1023_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2443_ _2125_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5231_ _0393_ net227 clknet_leaf_84_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5162_ _0324_ net206 clknet_leaf_88_clk net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_233_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2918__I Control_unit2.instr_stage2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4113_ _1611_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5093_ _0255_ net164 clknet_leaf_100_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_238_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _1453_ _1558_ _1564_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_237_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3661__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3749__I _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2653__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4946_ _0108_ net281 clknet_leaf_31_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_205_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__A1 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4877_ Control_unit1.instr_stage1\[12\] net147 clknet_leaf_13_clk Control_unit2.instr_stage2\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3828_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4875__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3484__I _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3759_ _1315_ _1366_ _1371_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4677__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4905__RN net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4429__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3659__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3394__I _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2391__A2 Control_unit2.instr_decoder2.A\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5149__RN net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__CLK clknet_leaf_66_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3891__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5180__CLK clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout175_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3643__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4800_ _0002_ net118 clknet_leaf_12_clk net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout342_I net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2992_ _0812_ _0813_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_222_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4731_ _1068_ _1414_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _1882_ _1987_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3159__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3613_ _1130_ _1259_ _1263_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4593_ _1920_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5388__RN net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3544_ _1163_ _1211_ _1217_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3475_ _1163_ _1154_ _1164_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5214_ _0376_ net224 clknet_leaf_80_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2426_ net37 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_213_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout88_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3331__A1 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5145_ _0307_ net207 clknet_leaf_87_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_245_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3882__A2 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5076_ _0238_ net180 clknet_leaf_104_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4027_ _1485_ _1550_ _1553_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_246_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4929_ _0091_ net266 clknet_leaf_27_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_200_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__RN net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3147__C _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3570__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3942__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output69_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3322__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5303__RN net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3389__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4050__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4013__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3260_ _0822_ _1000_ _1012_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3313__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3191_ _0832_ _0956_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_223_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2975_ _0795_ _0796_ _0800_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4041__A2 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4714_ _0998_ _2019_ _2021_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5076__CLK clknet_leaf_104_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4645_ _0933_ _1226_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5166__D _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4576_ _1885_ _1931_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _1138_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4913__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3458_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2409_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3389_ _1043_ _1100_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _0290_ net168 clknet_leaf_93_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input20_I read_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4593__I _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3068__B1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _0221_ net99 clknet_leaf_110_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3002__I _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4032__A2 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3138__A4 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3543__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3672__I _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4099__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4271__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5099__CLK clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2760_ Control_unit2.instr_decoder2.A\[1\] _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout138_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2585__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2691_ _2364_ _2371_ _2372_ _2373_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout305_I net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4430_ _1802_ _1825_ _1830_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4936__CLK clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3534__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__I _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4361_ _1733_ _1778_ _1786_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3312_ _0996_ _1049_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4292_ _1644_ _1729_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3243_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3837__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3174_ _2277_ _0943_ _0947_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2926__I Control_unit2.instr_stage2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_235_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4262__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4014__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2958_ _0786_ _0783_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2889_ _0706_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4628_ _1890_ _1965_ _1967_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3492__I _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4559_ _1864_ _1918_ _1922_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4809__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4253__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3667__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2571__I _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3064__I0 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4959__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4498__I _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_71_clk_I clknet_4_11_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput50 net50 instr_mem_addr[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput61 net61 write_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_218_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput72 net72 write_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3819__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2746__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4244__A2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3930_ _1343_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout255_I net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3861_ _1418_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_24_clk_I clknet_4_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2812_ Stack_pointer.SP\[6\] _0657_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3792_ _1360_ _1391_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2743_ _2206_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_203_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _2355_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_39_clk_I clknet_4_13_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5114__CLK clknet_leaf_88_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4413_ _1738_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5393_ _0555_ net118 clknet_leaf_6_clk net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ _1347_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout306 net308 net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout317 net319 net317 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2730__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout328 net352 net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout339 net351 net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_154_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4275_ _1630_ _1718_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5264__CLK clknet_leaf_77_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3226_ _0795_ _0982_ _0985_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_246_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4483__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3157_ _0934_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2494__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3088_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4786__A3 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3487__I _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2549__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_111_clk clknet_4_0_0_clk clknet_leaf_111_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4111__I _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output51_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2566__I _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2485__A1 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_clk clknet_4_9_0_clk clknet_leaf_102_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_220_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2390_ Arithmetic_Logic_Unit.op _2085_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3860__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4060_ _1473_ _1571_ _1574_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3011_ _0782_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4962_ _0124_ net267 clknet_leaf_27_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3913_ _1473_ _1469_ _1475_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3976__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4893_ net5 net146 clknet_leaf_15_clk Control_unit1.instr_stage1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2425__B _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3100__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3844_ _1308_ _1425_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_225_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3775_ _1336_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2726_ _2133_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_199_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2657_ _2317_ _2300_ _2326_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5174__D _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5376_ _0538_ net324 clknet_leaf_52_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2588_ _2276_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout103 net109 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout114 net117 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ net20 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout125 net126 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3770__I _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout136 net140 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout147 net151 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout158 net159 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4258_ _1606_ _1705_ _1710_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout169 net172 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_25_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3209_ _0962_ _0969_ _0972_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _1630_ _1664_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4106__I _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3010__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3680__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4447__A2 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout120_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4383__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ _1227_ _0881_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2511_ _2197_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_196_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3491_ _1174_ _1169_ _1177_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5230_ _0392_ net224 clknet_leaf_84_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2442_ _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_143_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4686__A2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5161_ _0323_ net207 clknet_leaf_88_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2697__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4112_ _1587_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5092_ _0254_ net161 clknet_leaf_103_clk net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4438__A2 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _1505_ _1560_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5302__CLK clknet_leaf_65_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _0107_ net281 clknet_leaf_31_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2621__A1 Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4876_ Control_unit1.instr_stage1\[11\] net147 clknet_leaf_13_clk Control_unit2.instr_stage2\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_221_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3827_ _0964_ _1414_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_197_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3758_ _1316_ _1367_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2924__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2709_ _0564_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3689_ _1315_ _1302_ _1317_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_238_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5359_ _0521_ net323 clknet_leaf_53_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_5905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3005__I _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__A2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2612__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__RN net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3675__I _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__A3 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5325__CLK clknet_leaf_59_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_234_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout168_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2991_ _0782_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ _1027_ _2025_ _2030_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_226_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4832__RN net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4661_ _1929_ _1986_ _1988_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3585__I _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3612_ _1196_ _1261_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4592_ _1917_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3543_ _1216_ _1212_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_196_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3474_ _1058_ _1157_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5213_ _0375_ net214 clknet_leaf_82_clk net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2425_ _2083_ _2118_ _2119_ _2101_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_237_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3331__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5144_ _0306_ net169 clknet_leaf_93_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4899__RN net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _0237_ net99 clknet_leaf_110_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_229_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4026_ _1486_ _1551_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3095__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_91_clk clknet_4_10_0_clk clknet_leaf_91_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_225_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4595__A1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _0090_ net343 clknet_leaf_46_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_212_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4823__RN net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ Stack_pointer.SP_next\[3\] net122 clknet_leaf_9_clk Stack_pointer.SP\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5348__CLK clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3322__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2833__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_82_clk clknet_4_11_0_clk clknet_leaf_82_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5067__RN net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3190_ _0571_ _0955_ _0957_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout285_I net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2824__A1 Control_unit1.instr_decoder1.A\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_73_clk clknet_4_14_0_clk clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_235_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4577__A1 _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5058__RN net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2974_ _0798_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_222_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__RN net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4713_ _0811_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4329__A1 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4644_ _1913_ _1971_ _1976_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4575_ _1881_ _1930_ _1933_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3552__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3526_ _1192_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3457_ net31 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2408_ _2101_ _2102_ _2093_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3388_ _0974_ _1098_ _1102_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5127_ _0289_ net167 clknet_leaf_95_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3068__A1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ _0220_ net99 clknet_leaf_110_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_input13_I instr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3068__B2 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4009_ _1462_ _1538_ _1542_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2815__A1 Stack_pointer.SP\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64_clk clknet_4_12_0_clk clknet_leaf_64_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4568__A1 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5020__CLK clknet_leaf_73_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3240__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5170__CLK clknet_leaf_113_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4740__A1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2569__I _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4888__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5288__RN net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_clk clknet_4_14_0_clk clknet_leaf_55_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4559__A1 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3782__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2690_ _2307_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_223_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout200_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__RN net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1785_ _1781_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3311_ _0991_ _1048_ _1052_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _1296_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3242_ _2321_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3298__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I instr[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_230_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3173_ _0805_ _0944_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_239_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__RN net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2648__I1 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_clk clknet_4_15_0_clk clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5043__CLK clknet_leaf_108_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2957_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5193__CLK clknet_leaf_94_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2888_ _0724_ _0725_ _0715_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_202_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4627_ _1892_ _1966_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3773__I _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5203__RN net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4558_ _1919_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3509_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4489_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4109__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_233_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_37_clk clknet_4_13_0_clk clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3213__A1 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3064__I1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4779__I _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4713__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput40 net40 data_mem_addr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput51 net76 instr_mem_addr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput62 net62 write_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_155_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput73 net73 write_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_28_clk clknet_4_3_0_clk clknet_leaf_28_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout150_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ _1416_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout248_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4903__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2811_ Stack_pointer.SP\[6\] _0657_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3791_ _1294_ _1389_ _1393_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2742_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[0\].i2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2673_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3 _2305_ _2356_ _2307_ _2357_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4412_ _1813_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4704__A1 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ _0554_ net325 clknet_leaf_52_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_201_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4343_ _1770_ _1763_ _1772_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout307 net308 net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_193_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout318 net320 net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout329 net332 net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4274_ _1626_ _1717_ _1720_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3225_ _0983_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3156_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_19_clk clknet_4_4_0_clk clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3087_ _0879_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3989_ _1528_ _1226_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3746__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3008__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5089__CLK clknet_leaf_109_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_246_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_246_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2582__I Arithmetic_Logic_Unit.ALU_001.Y_CY\[7\].i3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A2 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4302__I _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout198_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3010_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _0123_ net267 clknet_leaf_27_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2492__I _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3912_ _1474_ _1471_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4892_ net4 net125 clknet_leaf_10_clk Control_unit1.instr_stage1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_220_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3843_ _1365_ _1424_ _1426_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_225_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3774_ _1355_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _0572_ _0580_ _0582_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_88_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_clk clknet_4_5_0_clk clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2656_ _2249_ _2340_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5231__CLK clknet_leaf_84_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2587_ _2257_ _2270_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5375_ _0537_ net324 clknet_leaf_52_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout104 net107 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout115 net117 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4326_ _1758_ _1751_ _1759_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout126 net127 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_232_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout137 net140 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout148 net150 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5381__CLK clknet_leaf_28_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout159 net160 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4257_ _1607_ _1706_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4949__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3208_ _0781_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4188_ _1626_ _1663_ _1666_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_227_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3664__A1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3139_ _0599_ _0919_ _0865_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_70_clk_I clknet_4_9_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3498__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3719__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_85_clk_I clknet_4_10_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4122__I _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_clk_I clknet_4_13_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5254__CLK clknet_leaf_104_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4383__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2510_ _2198_ _2182_ _2201_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3490_ _1176_ _1172_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2441_ _2093_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5160_ _0322_ net169 clknet_leaf_93_clk net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2697__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4111_ _1155_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5091_ _0253_ net101 clknet_leaf_110_clk net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4042_ _1451_ _1558_ _1563_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_231_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3646__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4207__I _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3111__I _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4944_ _0106_ net342 clknet_leaf_46_clk net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4875_ Control_unit1.instr_stage1\[10\] net129 clknet_leaf_3_clk Control_unit2.instr_stage2\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_127_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2950__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3826_ _1228_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3757_ _1311_ _1366_ _1370_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2708_ _2160_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3688_ _1316_ _1304_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2639_ _2124_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[10\].i0 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5358_ _0520_ net321 clknet_leaf_51_clk net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4309_ _1744_ _1737_ _1746_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5289_ _0451_ net231 clknet_leaf_71_clk net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3637__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__CLK clknet_leaf_95_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4062__A1 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5277__CLK clknet_leaf_72_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2612__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3956__I _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3691__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3876__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2990_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2603__A2 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout230_I net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _1878_ _1987_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout328_I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3611_ _1123_ _1259_ _1262_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_200_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4591_ _1942_ _1936_ _1943_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3542_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3473_ _1008_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2424_ _2079_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5212_ _0374_ net175 clknet_leaf_91_clk net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5143_ _0305_ net167 clknet_leaf_95_clk net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _0236_ net99 clknet_leaf_109_clk net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4025_ _1480_ _1550_ _1552_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3095__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4292__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4927_ _0089_ net343 clknet_leaf_45_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4595__A2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4858_ Stack_pointer.SP_next\[2\] net116 clknet_leaf_9_clk Stack_pointer.SP\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_240_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3809_ _1319_ _1402_ _1404_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4347__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4789_ _2068_ _2070_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4400__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3858__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2530__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3686__I _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2590__I _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2597__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4338__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4310__I _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout180_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout278_I net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2973_ _0782_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3596__I _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4712_ _2007_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ _1914_ _1972_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4574_ _1882_ _1931_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3525_ _1188_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3456_ _0994_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2407_ _2081_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3387_ _1041_ _1100_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5126_ _0288_ net167 clknet_leaf_95_clk net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ _0219_ net180 clknet_leaf_103_clk net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4265__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4008_ _1463_ _1539_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4568__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5315__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output74_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2503__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4559__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4799__RN net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3310_ _0992_ _1049_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _1731_ _1727_ _1732_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4971__RN net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3241_ _0995_ _0982_ _0997_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4832__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3172_ _2256_ _0943_ _0946_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4247__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4982__CLK clknet_leaf_64_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5338__CLK clknet_leaf_62_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2956_ net25 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2887_ net79 _0723_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_176_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4626_ _1953_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4557_ _1920_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3508_ _1187_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4488_ _1865_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3439_ _1134_ _1126_ _1135_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _0271_ net163 clknet_leaf_100_clk net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_246_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4125__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4855__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput41 net41 data_mem_addr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput52 net52 instr_mem_addr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_194_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput63 net63 write_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput74 net74 write_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3204__I _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4035__I _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2810_ _0638_ _0640_ _0658_ _0660_ Stack_pointer.SP_next\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3790_ _1358_ _1391_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2741_ _0597_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3874__I _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout310_I net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _2124_ Arithmetic_Logic_Unit.ALU_001.Y_CY\[11\].i3 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _1811_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5391_ _0553_ net325 clknet_leaf_52_clk net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2715__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5197__RN net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4342_ _1771_ _1765_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout308 net314 net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout319 net320 net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4273_ _1627_ _1718_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5010__CLK clknet_leaf_107_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3224_ _0970_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

