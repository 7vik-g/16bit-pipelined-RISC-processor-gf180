magic
tech gf180mcuC
magscale 1 5
timestamp 1670490271
<< obsm1 >>
rect 672 855 99288 99553
<< metal2 >>
rect 7112 99600 7168 100000
rect 7448 99600 7504 100000
rect 7784 99600 7840 100000
rect 8120 99600 8176 100000
rect 8456 99600 8512 100000
rect 8792 99600 8848 100000
rect 9128 99600 9184 100000
rect 9464 99600 9520 100000
rect 9800 99600 9856 100000
rect 10136 99600 10192 100000
rect 10472 99600 10528 100000
rect 10808 99600 10864 100000
rect 11144 99600 11200 100000
rect 11480 99600 11536 100000
rect 11816 99600 11872 100000
rect 12152 99600 12208 100000
rect 12488 99600 12544 100000
rect 12824 99600 12880 100000
rect 13160 99600 13216 100000
rect 13496 99600 13552 100000
rect 13832 99600 13888 100000
rect 14168 99600 14224 100000
rect 14504 99600 14560 100000
rect 14840 99600 14896 100000
rect 15176 99600 15232 100000
rect 15512 99600 15568 100000
rect 15848 99600 15904 100000
rect 16184 99600 16240 100000
rect 16520 99600 16576 100000
rect 16856 99600 16912 100000
rect 17192 99600 17248 100000
rect 17528 99600 17584 100000
rect 17864 99600 17920 100000
rect 18200 99600 18256 100000
rect 18536 99600 18592 100000
rect 18872 99600 18928 100000
rect 19208 99600 19264 100000
rect 19544 99600 19600 100000
rect 19880 99600 19936 100000
rect 20216 99600 20272 100000
rect 20552 99600 20608 100000
rect 20888 99600 20944 100000
rect 21224 99600 21280 100000
rect 21560 99600 21616 100000
rect 21896 99600 21952 100000
rect 22232 99600 22288 100000
rect 22568 99600 22624 100000
rect 22904 99600 22960 100000
rect 23240 99600 23296 100000
rect 23576 99600 23632 100000
rect 23912 99600 23968 100000
rect 24248 99600 24304 100000
rect 24584 99600 24640 100000
rect 24920 99600 24976 100000
rect 25256 99600 25312 100000
rect 25592 99600 25648 100000
rect 25928 99600 25984 100000
rect 26264 99600 26320 100000
rect 26600 99600 26656 100000
rect 26936 99600 26992 100000
rect 27272 99600 27328 100000
rect 27608 99600 27664 100000
rect 27944 99600 28000 100000
rect 28280 99600 28336 100000
rect 28616 99600 28672 100000
rect 28952 99600 29008 100000
rect 29288 99600 29344 100000
rect 29624 99600 29680 100000
rect 29960 99600 30016 100000
rect 30296 99600 30352 100000
rect 30632 99600 30688 100000
rect 30968 99600 31024 100000
rect 31304 99600 31360 100000
rect 31640 99600 31696 100000
rect 31976 99600 32032 100000
rect 32312 99600 32368 100000
rect 32648 99600 32704 100000
rect 32984 99600 33040 100000
rect 33320 99600 33376 100000
rect 33656 99600 33712 100000
rect 33992 99600 34048 100000
rect 34328 99600 34384 100000
rect 34664 99600 34720 100000
rect 35000 99600 35056 100000
rect 35336 99600 35392 100000
rect 35672 99600 35728 100000
rect 36008 99600 36064 100000
rect 36344 99600 36400 100000
rect 36680 99600 36736 100000
rect 37016 99600 37072 100000
rect 37352 99600 37408 100000
rect 37688 99600 37744 100000
rect 38024 99600 38080 100000
rect 38360 99600 38416 100000
rect 38696 99600 38752 100000
rect 39032 99600 39088 100000
rect 39368 99600 39424 100000
rect 39704 99600 39760 100000
rect 40040 99600 40096 100000
rect 40376 99600 40432 100000
rect 40712 99600 40768 100000
rect 41048 99600 41104 100000
rect 41384 99600 41440 100000
rect 41720 99600 41776 100000
rect 42056 99600 42112 100000
rect 42392 99600 42448 100000
rect 42728 99600 42784 100000
rect 43064 99600 43120 100000
rect 43400 99600 43456 100000
rect 43736 99600 43792 100000
rect 44072 99600 44128 100000
rect 44408 99600 44464 100000
rect 44744 99600 44800 100000
rect 45080 99600 45136 100000
rect 45416 99600 45472 100000
rect 45752 99600 45808 100000
rect 46088 99600 46144 100000
rect 46424 99600 46480 100000
rect 46760 99600 46816 100000
rect 47096 99600 47152 100000
rect 47432 99600 47488 100000
rect 47768 99600 47824 100000
rect 48104 99600 48160 100000
rect 48440 99600 48496 100000
rect 48776 99600 48832 100000
rect 49112 99600 49168 100000
rect 49448 99600 49504 100000
rect 49784 99600 49840 100000
rect 50120 99600 50176 100000
rect 50456 99600 50512 100000
rect 50792 99600 50848 100000
rect 51128 99600 51184 100000
rect 51464 99600 51520 100000
rect 51800 99600 51856 100000
rect 52136 99600 52192 100000
rect 52472 99600 52528 100000
rect 52808 99600 52864 100000
rect 53144 99600 53200 100000
rect 53480 99600 53536 100000
rect 53816 99600 53872 100000
rect 54152 99600 54208 100000
rect 54488 99600 54544 100000
rect 54824 99600 54880 100000
rect 55160 99600 55216 100000
rect 55496 99600 55552 100000
rect 55832 99600 55888 100000
rect 56168 99600 56224 100000
rect 56504 99600 56560 100000
rect 56840 99600 56896 100000
rect 57176 99600 57232 100000
rect 57512 99600 57568 100000
rect 57848 99600 57904 100000
rect 58184 99600 58240 100000
rect 58520 99600 58576 100000
rect 58856 99600 58912 100000
rect 59192 99600 59248 100000
rect 59528 99600 59584 100000
rect 59864 99600 59920 100000
rect 60200 99600 60256 100000
rect 60536 99600 60592 100000
rect 60872 99600 60928 100000
rect 61208 99600 61264 100000
rect 61544 99600 61600 100000
rect 61880 99600 61936 100000
rect 62216 99600 62272 100000
rect 62552 99600 62608 100000
rect 62888 99600 62944 100000
rect 63224 99600 63280 100000
rect 63560 99600 63616 100000
rect 63896 99600 63952 100000
rect 64232 99600 64288 100000
rect 64568 99600 64624 100000
rect 64904 99600 64960 100000
rect 65240 99600 65296 100000
rect 65576 99600 65632 100000
rect 65912 99600 65968 100000
rect 66248 99600 66304 100000
rect 66584 99600 66640 100000
rect 66920 99600 66976 100000
rect 67256 99600 67312 100000
rect 67592 99600 67648 100000
rect 67928 99600 67984 100000
rect 68264 99600 68320 100000
rect 68600 99600 68656 100000
rect 68936 99600 68992 100000
rect 69272 99600 69328 100000
rect 69608 99600 69664 100000
rect 69944 99600 70000 100000
rect 70280 99600 70336 100000
rect 70616 99600 70672 100000
rect 70952 99600 71008 100000
rect 71288 99600 71344 100000
rect 71624 99600 71680 100000
rect 71960 99600 72016 100000
rect 72296 99600 72352 100000
rect 72632 99600 72688 100000
rect 72968 99600 73024 100000
rect 73304 99600 73360 100000
rect 73640 99600 73696 100000
rect 73976 99600 74032 100000
rect 74312 99600 74368 100000
rect 74648 99600 74704 100000
rect 74984 99600 75040 100000
rect 75320 99600 75376 100000
rect 75656 99600 75712 100000
rect 75992 99600 76048 100000
rect 76328 99600 76384 100000
rect 76664 99600 76720 100000
rect 77000 99600 77056 100000
rect 77336 99600 77392 100000
rect 77672 99600 77728 100000
rect 78008 99600 78064 100000
rect 78344 99600 78400 100000
rect 78680 99600 78736 100000
rect 79016 99600 79072 100000
rect 79352 99600 79408 100000
rect 79688 99600 79744 100000
rect 80024 99600 80080 100000
rect 80360 99600 80416 100000
rect 80696 99600 80752 100000
rect 81032 99600 81088 100000
rect 81368 99600 81424 100000
rect 81704 99600 81760 100000
rect 82040 99600 82096 100000
rect 82376 99600 82432 100000
rect 82712 99600 82768 100000
rect 83048 99600 83104 100000
rect 83384 99600 83440 100000
rect 83720 99600 83776 100000
rect 84056 99600 84112 100000
rect 84392 99600 84448 100000
rect 84728 99600 84784 100000
rect 85064 99600 85120 100000
rect 85400 99600 85456 100000
rect 85736 99600 85792 100000
rect 86072 99600 86128 100000
rect 86408 99600 86464 100000
rect 86744 99600 86800 100000
rect 87080 99600 87136 100000
rect 87416 99600 87472 100000
rect 87752 99600 87808 100000
rect 88088 99600 88144 100000
rect 88424 99600 88480 100000
rect 88760 99600 88816 100000
rect 89096 99600 89152 100000
rect 89432 99600 89488 100000
rect 89768 99600 89824 100000
rect 90104 99600 90160 100000
rect 90440 99600 90496 100000
rect 90776 99600 90832 100000
rect 91112 99600 91168 100000
rect 91448 99600 91504 100000
rect 91784 99600 91840 100000
rect 92120 99600 92176 100000
rect 92456 99600 92512 100000
rect 92792 99600 92848 100000
rect 784 0 840 400
rect 1512 0 1568 400
rect 2240 0 2296 400
rect 2968 0 3024 400
rect 3696 0 3752 400
rect 4424 0 4480 400
rect 5152 0 5208 400
rect 5880 0 5936 400
rect 6608 0 6664 400
rect 7336 0 7392 400
rect 8064 0 8120 400
rect 8792 0 8848 400
rect 9520 0 9576 400
rect 10248 0 10304 400
rect 10976 0 11032 400
rect 11704 0 11760 400
rect 12432 0 12488 400
rect 13160 0 13216 400
rect 13888 0 13944 400
rect 14616 0 14672 400
rect 15344 0 15400 400
rect 16072 0 16128 400
rect 16800 0 16856 400
rect 17528 0 17584 400
rect 18256 0 18312 400
rect 18984 0 19040 400
rect 19712 0 19768 400
rect 20440 0 20496 400
rect 21168 0 21224 400
rect 21896 0 21952 400
rect 22624 0 22680 400
rect 23352 0 23408 400
rect 24080 0 24136 400
rect 24808 0 24864 400
rect 25536 0 25592 400
rect 26264 0 26320 400
rect 26992 0 27048 400
rect 27720 0 27776 400
rect 28448 0 28504 400
rect 29176 0 29232 400
rect 29904 0 29960 400
rect 30632 0 30688 400
rect 31360 0 31416 400
rect 32088 0 32144 400
rect 32816 0 32872 400
rect 33544 0 33600 400
rect 34272 0 34328 400
rect 35000 0 35056 400
rect 35728 0 35784 400
rect 36456 0 36512 400
rect 37184 0 37240 400
rect 37912 0 37968 400
rect 38640 0 38696 400
rect 39368 0 39424 400
rect 40096 0 40152 400
rect 40824 0 40880 400
rect 41552 0 41608 400
rect 42280 0 42336 400
rect 43008 0 43064 400
rect 43736 0 43792 400
rect 44464 0 44520 400
rect 45192 0 45248 400
rect 45920 0 45976 400
rect 46648 0 46704 400
rect 47376 0 47432 400
rect 48104 0 48160 400
rect 48832 0 48888 400
rect 49560 0 49616 400
rect 50288 0 50344 400
rect 51016 0 51072 400
rect 51744 0 51800 400
rect 52472 0 52528 400
rect 53200 0 53256 400
rect 53928 0 53984 400
rect 54656 0 54712 400
rect 55384 0 55440 400
rect 56112 0 56168 400
rect 56840 0 56896 400
rect 57568 0 57624 400
rect 58296 0 58352 400
rect 59024 0 59080 400
rect 59752 0 59808 400
rect 60480 0 60536 400
rect 61208 0 61264 400
rect 61936 0 61992 400
rect 62664 0 62720 400
rect 63392 0 63448 400
rect 64120 0 64176 400
rect 64848 0 64904 400
rect 65576 0 65632 400
rect 66304 0 66360 400
rect 67032 0 67088 400
rect 67760 0 67816 400
rect 68488 0 68544 400
rect 69216 0 69272 400
rect 69944 0 70000 400
rect 70672 0 70728 400
rect 71400 0 71456 400
rect 72128 0 72184 400
rect 72856 0 72912 400
rect 73584 0 73640 400
rect 74312 0 74368 400
rect 75040 0 75096 400
rect 75768 0 75824 400
rect 76496 0 76552 400
rect 77224 0 77280 400
rect 77952 0 78008 400
rect 78680 0 78736 400
rect 79408 0 79464 400
rect 80136 0 80192 400
rect 80864 0 80920 400
rect 81592 0 81648 400
rect 82320 0 82376 400
rect 83048 0 83104 400
rect 83776 0 83832 400
rect 84504 0 84560 400
rect 85232 0 85288 400
rect 85960 0 86016 400
rect 86688 0 86744 400
rect 87416 0 87472 400
rect 88144 0 88200 400
rect 88872 0 88928 400
rect 89600 0 89656 400
rect 90328 0 90384 400
rect 91056 0 91112 400
rect 91784 0 91840 400
rect 92512 0 92568 400
rect 93240 0 93296 400
rect 93968 0 94024 400
rect 94696 0 94752 400
rect 95424 0 95480 400
rect 96152 0 96208 400
rect 96880 0 96936 400
rect 97608 0 97664 400
rect 98336 0 98392 400
rect 99064 0 99120 400
<< obsm2 >>
rect 798 99570 7082 99951
rect 7198 99570 7418 99951
rect 7534 99570 7754 99951
rect 7870 99570 8090 99951
rect 8206 99570 8426 99951
rect 8542 99570 8762 99951
rect 8878 99570 9098 99951
rect 9214 99570 9434 99951
rect 9550 99570 9770 99951
rect 9886 99570 10106 99951
rect 10222 99570 10442 99951
rect 10558 99570 10778 99951
rect 10894 99570 11114 99951
rect 11230 99570 11450 99951
rect 11566 99570 11786 99951
rect 11902 99570 12122 99951
rect 12238 99570 12458 99951
rect 12574 99570 12794 99951
rect 12910 99570 13130 99951
rect 13246 99570 13466 99951
rect 13582 99570 13802 99951
rect 13918 99570 14138 99951
rect 14254 99570 14474 99951
rect 14590 99570 14810 99951
rect 14926 99570 15146 99951
rect 15262 99570 15482 99951
rect 15598 99570 15818 99951
rect 15934 99570 16154 99951
rect 16270 99570 16490 99951
rect 16606 99570 16826 99951
rect 16942 99570 17162 99951
rect 17278 99570 17498 99951
rect 17614 99570 17834 99951
rect 17950 99570 18170 99951
rect 18286 99570 18506 99951
rect 18622 99570 18842 99951
rect 18958 99570 19178 99951
rect 19294 99570 19514 99951
rect 19630 99570 19850 99951
rect 19966 99570 20186 99951
rect 20302 99570 20522 99951
rect 20638 99570 20858 99951
rect 20974 99570 21194 99951
rect 21310 99570 21530 99951
rect 21646 99570 21866 99951
rect 21982 99570 22202 99951
rect 22318 99570 22538 99951
rect 22654 99570 22874 99951
rect 22990 99570 23210 99951
rect 23326 99570 23546 99951
rect 23662 99570 23882 99951
rect 23998 99570 24218 99951
rect 24334 99570 24554 99951
rect 24670 99570 24890 99951
rect 25006 99570 25226 99951
rect 25342 99570 25562 99951
rect 25678 99570 25898 99951
rect 26014 99570 26234 99951
rect 26350 99570 26570 99951
rect 26686 99570 26906 99951
rect 27022 99570 27242 99951
rect 27358 99570 27578 99951
rect 27694 99570 27914 99951
rect 28030 99570 28250 99951
rect 28366 99570 28586 99951
rect 28702 99570 28922 99951
rect 29038 99570 29258 99951
rect 29374 99570 29594 99951
rect 29710 99570 29930 99951
rect 30046 99570 30266 99951
rect 30382 99570 30602 99951
rect 30718 99570 30938 99951
rect 31054 99570 31274 99951
rect 31390 99570 31610 99951
rect 31726 99570 31946 99951
rect 32062 99570 32282 99951
rect 32398 99570 32618 99951
rect 32734 99570 32954 99951
rect 33070 99570 33290 99951
rect 33406 99570 33626 99951
rect 33742 99570 33962 99951
rect 34078 99570 34298 99951
rect 34414 99570 34634 99951
rect 34750 99570 34970 99951
rect 35086 99570 35306 99951
rect 35422 99570 35642 99951
rect 35758 99570 35978 99951
rect 36094 99570 36314 99951
rect 36430 99570 36650 99951
rect 36766 99570 36986 99951
rect 37102 99570 37322 99951
rect 37438 99570 37658 99951
rect 37774 99570 37994 99951
rect 38110 99570 38330 99951
rect 38446 99570 38666 99951
rect 38782 99570 39002 99951
rect 39118 99570 39338 99951
rect 39454 99570 39674 99951
rect 39790 99570 40010 99951
rect 40126 99570 40346 99951
rect 40462 99570 40682 99951
rect 40798 99570 41018 99951
rect 41134 99570 41354 99951
rect 41470 99570 41690 99951
rect 41806 99570 42026 99951
rect 42142 99570 42362 99951
rect 42478 99570 42698 99951
rect 42814 99570 43034 99951
rect 43150 99570 43370 99951
rect 43486 99570 43706 99951
rect 43822 99570 44042 99951
rect 44158 99570 44378 99951
rect 44494 99570 44714 99951
rect 44830 99570 45050 99951
rect 45166 99570 45386 99951
rect 45502 99570 45722 99951
rect 45838 99570 46058 99951
rect 46174 99570 46394 99951
rect 46510 99570 46730 99951
rect 46846 99570 47066 99951
rect 47182 99570 47402 99951
rect 47518 99570 47738 99951
rect 47854 99570 48074 99951
rect 48190 99570 48410 99951
rect 48526 99570 48746 99951
rect 48862 99570 49082 99951
rect 49198 99570 49418 99951
rect 49534 99570 49754 99951
rect 49870 99570 50090 99951
rect 50206 99570 50426 99951
rect 50542 99570 50762 99951
rect 50878 99570 51098 99951
rect 51214 99570 51434 99951
rect 51550 99570 51770 99951
rect 51886 99570 52106 99951
rect 52222 99570 52442 99951
rect 52558 99570 52778 99951
rect 52894 99570 53114 99951
rect 53230 99570 53450 99951
rect 53566 99570 53786 99951
rect 53902 99570 54122 99951
rect 54238 99570 54458 99951
rect 54574 99570 54794 99951
rect 54910 99570 55130 99951
rect 55246 99570 55466 99951
rect 55582 99570 55802 99951
rect 55918 99570 56138 99951
rect 56254 99570 56474 99951
rect 56590 99570 56810 99951
rect 56926 99570 57146 99951
rect 57262 99570 57482 99951
rect 57598 99570 57818 99951
rect 57934 99570 58154 99951
rect 58270 99570 58490 99951
rect 58606 99570 58826 99951
rect 58942 99570 59162 99951
rect 59278 99570 59498 99951
rect 59614 99570 59834 99951
rect 59950 99570 60170 99951
rect 60286 99570 60506 99951
rect 60622 99570 60842 99951
rect 60958 99570 61178 99951
rect 61294 99570 61514 99951
rect 61630 99570 61850 99951
rect 61966 99570 62186 99951
rect 62302 99570 62522 99951
rect 62638 99570 62858 99951
rect 62974 99570 63194 99951
rect 63310 99570 63530 99951
rect 63646 99570 63866 99951
rect 63982 99570 64202 99951
rect 64318 99570 64538 99951
rect 64654 99570 64874 99951
rect 64990 99570 65210 99951
rect 65326 99570 65546 99951
rect 65662 99570 65882 99951
rect 65998 99570 66218 99951
rect 66334 99570 66554 99951
rect 66670 99570 66890 99951
rect 67006 99570 67226 99951
rect 67342 99570 67562 99951
rect 67678 99570 67898 99951
rect 68014 99570 68234 99951
rect 68350 99570 68570 99951
rect 68686 99570 68906 99951
rect 69022 99570 69242 99951
rect 69358 99570 69578 99951
rect 69694 99570 69914 99951
rect 70030 99570 70250 99951
rect 70366 99570 70586 99951
rect 70702 99570 70922 99951
rect 71038 99570 71258 99951
rect 71374 99570 71594 99951
rect 71710 99570 71930 99951
rect 72046 99570 72266 99951
rect 72382 99570 72602 99951
rect 72718 99570 72938 99951
rect 73054 99570 73274 99951
rect 73390 99570 73610 99951
rect 73726 99570 73946 99951
rect 74062 99570 74282 99951
rect 74398 99570 74618 99951
rect 74734 99570 74954 99951
rect 75070 99570 75290 99951
rect 75406 99570 75626 99951
rect 75742 99570 75962 99951
rect 76078 99570 76298 99951
rect 76414 99570 76634 99951
rect 76750 99570 76970 99951
rect 77086 99570 77306 99951
rect 77422 99570 77642 99951
rect 77758 99570 77978 99951
rect 78094 99570 78314 99951
rect 78430 99570 78650 99951
rect 78766 99570 78986 99951
rect 79102 99570 79322 99951
rect 79438 99570 79658 99951
rect 79774 99570 79994 99951
rect 80110 99570 80330 99951
rect 80446 99570 80666 99951
rect 80782 99570 81002 99951
rect 81118 99570 81338 99951
rect 81454 99570 81674 99951
rect 81790 99570 82010 99951
rect 82126 99570 82346 99951
rect 82462 99570 82682 99951
rect 82798 99570 83018 99951
rect 83134 99570 83354 99951
rect 83470 99570 83690 99951
rect 83806 99570 84026 99951
rect 84142 99570 84362 99951
rect 84478 99570 84698 99951
rect 84814 99570 85034 99951
rect 85150 99570 85370 99951
rect 85486 99570 85706 99951
rect 85822 99570 86042 99951
rect 86158 99570 86378 99951
rect 86494 99570 86714 99951
rect 86830 99570 87050 99951
rect 87166 99570 87386 99951
rect 87502 99570 87722 99951
rect 87838 99570 88058 99951
rect 88174 99570 88394 99951
rect 88510 99570 88730 99951
rect 88846 99570 89066 99951
rect 89182 99570 89402 99951
rect 89518 99570 89738 99951
rect 89854 99570 90074 99951
rect 90190 99570 90410 99951
rect 90526 99570 90746 99951
rect 90862 99570 91082 99951
rect 91198 99570 91418 99951
rect 91534 99570 91754 99951
rect 91870 99570 92090 99951
rect 92206 99570 92426 99951
rect 92542 99570 92762 99951
rect 92878 99570 99162 99951
rect 798 430 99162 99570
rect 870 400 1482 430
rect 1598 400 2210 430
rect 2326 400 2938 430
rect 3054 400 3666 430
rect 3782 400 4394 430
rect 4510 400 5122 430
rect 5238 400 5850 430
rect 5966 400 6578 430
rect 6694 400 7306 430
rect 7422 400 8034 430
rect 8150 400 8762 430
rect 8878 400 9490 430
rect 9606 400 10218 430
rect 10334 400 10946 430
rect 11062 400 11674 430
rect 11790 400 12402 430
rect 12518 400 13130 430
rect 13246 400 13858 430
rect 13974 400 14586 430
rect 14702 400 15314 430
rect 15430 400 16042 430
rect 16158 400 16770 430
rect 16886 400 17498 430
rect 17614 400 18226 430
rect 18342 400 18954 430
rect 19070 400 19682 430
rect 19798 400 20410 430
rect 20526 400 21138 430
rect 21254 400 21866 430
rect 21982 400 22594 430
rect 22710 400 23322 430
rect 23438 400 24050 430
rect 24166 400 24778 430
rect 24894 400 25506 430
rect 25622 400 26234 430
rect 26350 400 26962 430
rect 27078 400 27690 430
rect 27806 400 28418 430
rect 28534 400 29146 430
rect 29262 400 29874 430
rect 29990 400 30602 430
rect 30718 400 31330 430
rect 31446 400 32058 430
rect 32174 400 32786 430
rect 32902 400 33514 430
rect 33630 400 34242 430
rect 34358 400 34970 430
rect 35086 400 35698 430
rect 35814 400 36426 430
rect 36542 400 37154 430
rect 37270 400 37882 430
rect 37998 400 38610 430
rect 38726 400 39338 430
rect 39454 400 40066 430
rect 40182 400 40794 430
rect 40910 400 41522 430
rect 41638 400 42250 430
rect 42366 400 42978 430
rect 43094 400 43706 430
rect 43822 400 44434 430
rect 44550 400 45162 430
rect 45278 400 45890 430
rect 46006 400 46618 430
rect 46734 400 47346 430
rect 47462 400 48074 430
rect 48190 400 48802 430
rect 48918 400 49530 430
rect 49646 400 50258 430
rect 50374 400 50986 430
rect 51102 400 51714 430
rect 51830 400 52442 430
rect 52558 400 53170 430
rect 53286 400 53898 430
rect 54014 400 54626 430
rect 54742 400 55354 430
rect 55470 400 56082 430
rect 56198 400 56810 430
rect 56926 400 57538 430
rect 57654 400 58266 430
rect 58382 400 58994 430
rect 59110 400 59722 430
rect 59838 400 60450 430
rect 60566 400 61178 430
rect 61294 400 61906 430
rect 62022 400 62634 430
rect 62750 400 63362 430
rect 63478 400 64090 430
rect 64206 400 64818 430
rect 64934 400 65546 430
rect 65662 400 66274 430
rect 66390 400 67002 430
rect 67118 400 67730 430
rect 67846 400 68458 430
rect 68574 400 69186 430
rect 69302 400 69914 430
rect 70030 400 70642 430
rect 70758 400 71370 430
rect 71486 400 72098 430
rect 72214 400 72826 430
rect 72942 400 73554 430
rect 73670 400 74282 430
rect 74398 400 75010 430
rect 75126 400 75738 430
rect 75854 400 76466 430
rect 76582 400 77194 430
rect 77310 400 77922 430
rect 78038 400 78650 430
rect 78766 400 79378 430
rect 79494 400 80106 430
rect 80222 400 80834 430
rect 80950 400 81562 430
rect 81678 400 82290 430
rect 82406 400 83018 430
rect 83134 400 83746 430
rect 83862 400 84474 430
rect 84590 400 85202 430
rect 85318 400 85930 430
rect 86046 400 86658 430
rect 86774 400 87386 430
rect 87502 400 88114 430
rect 88230 400 88842 430
rect 88958 400 89570 430
rect 89686 400 90298 430
rect 90414 400 91026 430
rect 91142 400 91754 430
rect 91870 400 92482 430
rect 92598 400 93210 430
rect 93326 400 93938 430
rect 94054 400 94666 430
rect 94782 400 95394 430
rect 95510 400 96122 430
rect 96238 400 96850 430
rect 96966 400 97578 430
rect 97694 400 98306 430
rect 98422 400 99034 430
rect 99150 400 99162 430
<< obsm3 >>
rect 1073 854 99167 99946
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
rect 94384 1538 94544 98422
<< obsm4 >>
rect 42238 98452 67242 99895
rect 42238 2249 48274 98452
rect 48494 2249 55954 98452
rect 56174 2249 63634 98452
rect 63854 2249 67242 98452
<< labels >>
rlabel metal2 s 97608 0 97664 400 6 clk
port 1 nsew signal output
rlabel metal2 s 63896 99600 63952 100000 6 data_mem_addr[0]
port 2 nsew signal output
rlabel metal2 s 64904 99600 64960 100000 6 data_mem_addr[1]
port 3 nsew signal output
rlabel metal2 s 65912 99600 65968 100000 6 data_mem_addr[2]
port 4 nsew signal output
rlabel metal2 s 66920 99600 66976 100000 6 data_mem_addr[3]
port 5 nsew signal output
rlabel metal2 s 67928 99600 67984 100000 6 data_mem_addr[4]
port 6 nsew signal output
rlabel metal2 s 68936 99600 68992 100000 6 data_mem_addr[5]
port 7 nsew signal output
rlabel metal2 s 69944 99600 70000 100000 6 data_mem_addr[6]
port 8 nsew signal output
rlabel metal2 s 70952 99600 71008 100000 6 data_mem_addr[7]
port 9 nsew signal output
rlabel metal2 s 64232 99600 64288 100000 6 data_read_data[0]
port 10 nsew signal input
rlabel metal2 s 73304 99600 73360 100000 6 data_read_data[10]
port 11 nsew signal input
rlabel metal2 s 73976 99600 74032 100000 6 data_read_data[11]
port 12 nsew signal input
rlabel metal2 s 74648 99600 74704 100000 6 data_read_data[12]
port 13 nsew signal input
rlabel metal2 s 75320 99600 75376 100000 6 data_read_data[13]
port 14 nsew signal input
rlabel metal2 s 75992 99600 76048 100000 6 data_read_data[14]
port 15 nsew signal input
rlabel metal2 s 76664 99600 76720 100000 6 data_read_data[15]
port 16 nsew signal input
rlabel metal2 s 65240 99600 65296 100000 6 data_read_data[1]
port 17 nsew signal input
rlabel metal2 s 66248 99600 66304 100000 6 data_read_data[2]
port 18 nsew signal input
rlabel metal2 s 67256 99600 67312 100000 6 data_read_data[3]
port 19 nsew signal input
rlabel metal2 s 68264 99600 68320 100000 6 data_read_data[4]
port 20 nsew signal input
rlabel metal2 s 69272 99600 69328 100000 6 data_read_data[5]
port 21 nsew signal input
rlabel metal2 s 70280 99600 70336 100000 6 data_read_data[6]
port 22 nsew signal input
rlabel metal2 s 71288 99600 71344 100000 6 data_read_data[7]
port 23 nsew signal input
rlabel metal2 s 71960 99600 72016 100000 6 data_read_data[8]
port 24 nsew signal input
rlabel metal2 s 72632 99600 72688 100000 6 data_read_data[9]
port 25 nsew signal input
rlabel metal2 s 64568 99600 64624 100000 6 data_write_data[0]
port 26 nsew signal output
rlabel metal2 s 73640 99600 73696 100000 6 data_write_data[10]
port 27 nsew signal output
rlabel metal2 s 74312 99600 74368 100000 6 data_write_data[11]
port 28 nsew signal output
rlabel metal2 s 74984 99600 75040 100000 6 data_write_data[12]
port 29 nsew signal output
rlabel metal2 s 75656 99600 75712 100000 6 data_write_data[13]
port 30 nsew signal output
rlabel metal2 s 76328 99600 76384 100000 6 data_write_data[14]
port 31 nsew signal output
rlabel metal2 s 77000 99600 77056 100000 6 data_write_data[15]
port 32 nsew signal output
rlabel metal2 s 65576 99600 65632 100000 6 data_write_data[1]
port 33 nsew signal output
rlabel metal2 s 66584 99600 66640 100000 6 data_write_data[2]
port 34 nsew signal output
rlabel metal2 s 67592 99600 67648 100000 6 data_write_data[3]
port 35 nsew signal output
rlabel metal2 s 68600 99600 68656 100000 6 data_write_data[4]
port 36 nsew signal output
rlabel metal2 s 69608 99600 69664 100000 6 data_write_data[5]
port 37 nsew signal output
rlabel metal2 s 70616 99600 70672 100000 6 data_write_data[6]
port 38 nsew signal output
rlabel metal2 s 71624 99600 71680 100000 6 data_write_data[7]
port 39 nsew signal output
rlabel metal2 s 72296 99600 72352 100000 6 data_write_data[8]
port 40 nsew signal output
rlabel metal2 s 72968 99600 73024 100000 6 data_write_data[9]
port 41 nsew signal output
rlabel metal2 s 63560 99600 63616 100000 6 dataw_en
port 42 nsew signal output
rlabel metal2 s 92792 99600 92848 100000 6 hlt
port 43 nsew signal input
rlabel metal2 s 77672 99600 77728 100000 6 instr[0]
port 44 nsew signal input
rlabel metal2 s 87752 99600 87808 100000 6 instr[10]
port 45 nsew signal input
rlabel metal2 s 88760 99600 88816 100000 6 instr[11]
port 46 nsew signal input
rlabel metal2 s 89768 99600 89824 100000 6 instr[12]
port 47 nsew signal input
rlabel metal2 s 90776 99600 90832 100000 6 instr[13]
port 48 nsew signal input
rlabel metal2 s 91448 99600 91504 100000 6 instr[14]
port 49 nsew signal input
rlabel metal2 s 92120 99600 92176 100000 6 instr[15]
port 50 nsew signal input
rlabel metal2 s 78680 99600 78736 100000 6 instr[1]
port 51 nsew signal input
rlabel metal2 s 79688 99600 79744 100000 6 instr[2]
port 52 nsew signal input
rlabel metal2 s 80696 99600 80752 100000 6 instr[3]
port 53 nsew signal input
rlabel metal2 s 81704 99600 81760 100000 6 instr[4]
port 54 nsew signal input
rlabel metal2 s 82712 99600 82768 100000 6 instr[5]
port 55 nsew signal input
rlabel metal2 s 83720 99600 83776 100000 6 instr[6]
port 56 nsew signal input
rlabel metal2 s 84728 99600 84784 100000 6 instr[7]
port 57 nsew signal input
rlabel metal2 s 85736 99600 85792 100000 6 instr[8]
port 58 nsew signal input
rlabel metal2 s 86744 99600 86800 100000 6 instr[9]
port 59 nsew signal input
rlabel metal2 s 78008 99600 78064 100000 6 instr_mem_addr[0]
port 60 nsew signal output
rlabel metal2 s 88088 99600 88144 100000 6 instr_mem_addr[10]
port 61 nsew signal output
rlabel metal2 s 89096 99600 89152 100000 6 instr_mem_addr[11]
port 62 nsew signal output
rlabel metal2 s 90104 99600 90160 100000 6 instr_mem_addr[12]
port 63 nsew signal output
rlabel metal2 s 79016 99600 79072 100000 6 instr_mem_addr[1]
port 64 nsew signal output
rlabel metal2 s 80024 99600 80080 100000 6 instr_mem_addr[2]
port 65 nsew signal output
rlabel metal2 s 81032 99600 81088 100000 6 instr_mem_addr[3]
port 66 nsew signal output
rlabel metal2 s 82040 99600 82096 100000 6 instr_mem_addr[4]
port 67 nsew signal output
rlabel metal2 s 83048 99600 83104 100000 6 instr_mem_addr[5]
port 68 nsew signal output
rlabel metal2 s 84056 99600 84112 100000 6 instr_mem_addr[6]
port 69 nsew signal output
rlabel metal2 s 85064 99600 85120 100000 6 instr_mem_addr[7]
port 70 nsew signal output
rlabel metal2 s 86072 99600 86128 100000 6 instr_mem_addr[8]
port 71 nsew signal output
rlabel metal2 s 87080 99600 87136 100000 6 instr_mem_addr[9]
port 72 nsew signal output
rlabel metal2 s 78344 99600 78400 100000 6 instr_write_data[0]
port 73 nsew signal output
rlabel metal2 s 88424 99600 88480 100000 6 instr_write_data[10]
port 74 nsew signal output
rlabel metal2 s 89432 99600 89488 100000 6 instr_write_data[11]
port 75 nsew signal output
rlabel metal2 s 90440 99600 90496 100000 6 instr_write_data[12]
port 76 nsew signal output
rlabel metal2 s 91112 99600 91168 100000 6 instr_write_data[13]
port 77 nsew signal output
rlabel metal2 s 91784 99600 91840 100000 6 instr_write_data[14]
port 78 nsew signal output
rlabel metal2 s 92456 99600 92512 100000 6 instr_write_data[15]
port 79 nsew signal output
rlabel metal2 s 79352 99600 79408 100000 6 instr_write_data[1]
port 80 nsew signal output
rlabel metal2 s 80360 99600 80416 100000 6 instr_write_data[2]
port 81 nsew signal output
rlabel metal2 s 81368 99600 81424 100000 6 instr_write_data[3]
port 82 nsew signal output
rlabel metal2 s 82376 99600 82432 100000 6 instr_write_data[4]
port 83 nsew signal output
rlabel metal2 s 83384 99600 83440 100000 6 instr_write_data[5]
port 84 nsew signal output
rlabel metal2 s 84392 99600 84448 100000 6 instr_write_data[6]
port 85 nsew signal output
rlabel metal2 s 85400 99600 85456 100000 6 instr_write_data[7]
port 86 nsew signal output
rlabel metal2 s 86408 99600 86464 100000 6 instr_write_data[8]
port 87 nsew signal output
rlabel metal2 s 87416 99600 87472 100000 6 instr_write_data[9]
port 88 nsew signal output
rlabel metal2 s 77336 99600 77392 100000 6 instrw_en
port 89 nsew signal output
rlabel metal2 s 7112 99600 7168 100000 6 io_in[0]
port 90 nsew signal input
rlabel metal2 s 17192 99600 17248 100000 6 io_in[10]
port 91 nsew signal input
rlabel metal2 s 18200 99600 18256 100000 6 io_in[11]
port 92 nsew signal input
rlabel metal2 s 19208 99600 19264 100000 6 io_in[12]
port 93 nsew signal input
rlabel metal2 s 20216 99600 20272 100000 6 io_in[13]
port 94 nsew signal input
rlabel metal2 s 21224 99600 21280 100000 6 io_in[14]
port 95 nsew signal input
rlabel metal2 s 22232 99600 22288 100000 6 io_in[15]
port 96 nsew signal input
rlabel metal2 s 23240 99600 23296 100000 6 io_in[16]
port 97 nsew signal input
rlabel metal2 s 24248 99600 24304 100000 6 io_in[17]
port 98 nsew signal input
rlabel metal2 s 25256 99600 25312 100000 6 io_in[18]
port 99 nsew signal input
rlabel metal2 s 26264 99600 26320 100000 6 io_in[19]
port 100 nsew signal input
rlabel metal2 s 8120 99600 8176 100000 6 io_in[1]
port 101 nsew signal input
rlabel metal2 s 27272 99600 27328 100000 6 io_in[20]
port 102 nsew signal input
rlabel metal2 s 28280 99600 28336 100000 6 io_in[21]
port 103 nsew signal input
rlabel metal2 s 29288 99600 29344 100000 6 io_in[22]
port 104 nsew signal input
rlabel metal2 s 30296 99600 30352 100000 6 io_in[23]
port 105 nsew signal input
rlabel metal2 s 31304 99600 31360 100000 6 io_in[24]
port 106 nsew signal input
rlabel metal2 s 32312 99600 32368 100000 6 io_in[25]
port 107 nsew signal input
rlabel metal2 s 33320 99600 33376 100000 6 io_in[26]
port 108 nsew signal input
rlabel metal2 s 34328 99600 34384 100000 6 io_in[27]
port 109 nsew signal input
rlabel metal2 s 35336 99600 35392 100000 6 io_in[28]
port 110 nsew signal input
rlabel metal2 s 36344 99600 36400 100000 6 io_in[29]
port 111 nsew signal input
rlabel metal2 s 9128 99600 9184 100000 6 io_in[2]
port 112 nsew signal input
rlabel metal2 s 37352 99600 37408 100000 6 io_in[30]
port 113 nsew signal input
rlabel metal2 s 38360 99600 38416 100000 6 io_in[31]
port 114 nsew signal input
rlabel metal2 s 39368 99600 39424 100000 6 io_in[32]
port 115 nsew signal input
rlabel metal2 s 40376 99600 40432 100000 6 io_in[33]
port 116 nsew signal input
rlabel metal2 s 41384 99600 41440 100000 6 io_in[34]
port 117 nsew signal input
rlabel metal2 s 42392 99600 42448 100000 6 io_in[35]
port 118 nsew signal input
rlabel metal2 s 43400 99600 43456 100000 6 io_in[36]
port 119 nsew signal input
rlabel metal2 s 44408 99600 44464 100000 6 io_in[37]
port 120 nsew signal input
rlabel metal2 s 10136 99600 10192 100000 6 io_in[3]
port 121 nsew signal input
rlabel metal2 s 11144 99600 11200 100000 6 io_in[4]
port 122 nsew signal input
rlabel metal2 s 12152 99600 12208 100000 6 io_in[5]
port 123 nsew signal input
rlabel metal2 s 13160 99600 13216 100000 6 io_in[6]
port 124 nsew signal input
rlabel metal2 s 14168 99600 14224 100000 6 io_in[7]
port 125 nsew signal input
rlabel metal2 s 15176 99600 15232 100000 6 io_in[8]
port 126 nsew signal input
rlabel metal2 s 16184 99600 16240 100000 6 io_in[9]
port 127 nsew signal input
rlabel metal2 s 7448 99600 7504 100000 6 io_oeb[0]
port 128 nsew signal output
rlabel metal2 s 17528 99600 17584 100000 6 io_oeb[10]
port 129 nsew signal output
rlabel metal2 s 18536 99600 18592 100000 6 io_oeb[11]
port 130 nsew signal output
rlabel metal2 s 19544 99600 19600 100000 6 io_oeb[12]
port 131 nsew signal output
rlabel metal2 s 20552 99600 20608 100000 6 io_oeb[13]
port 132 nsew signal output
rlabel metal2 s 21560 99600 21616 100000 6 io_oeb[14]
port 133 nsew signal output
rlabel metal2 s 22568 99600 22624 100000 6 io_oeb[15]
port 134 nsew signal output
rlabel metal2 s 23576 99600 23632 100000 6 io_oeb[16]
port 135 nsew signal output
rlabel metal2 s 24584 99600 24640 100000 6 io_oeb[17]
port 136 nsew signal output
rlabel metal2 s 25592 99600 25648 100000 6 io_oeb[18]
port 137 nsew signal output
rlabel metal2 s 26600 99600 26656 100000 6 io_oeb[19]
port 138 nsew signal output
rlabel metal2 s 8456 99600 8512 100000 6 io_oeb[1]
port 139 nsew signal output
rlabel metal2 s 27608 99600 27664 100000 6 io_oeb[20]
port 140 nsew signal output
rlabel metal2 s 28616 99600 28672 100000 6 io_oeb[21]
port 141 nsew signal output
rlabel metal2 s 29624 99600 29680 100000 6 io_oeb[22]
port 142 nsew signal output
rlabel metal2 s 30632 99600 30688 100000 6 io_oeb[23]
port 143 nsew signal output
rlabel metal2 s 31640 99600 31696 100000 6 io_oeb[24]
port 144 nsew signal output
rlabel metal2 s 32648 99600 32704 100000 6 io_oeb[25]
port 145 nsew signal output
rlabel metal2 s 33656 99600 33712 100000 6 io_oeb[26]
port 146 nsew signal output
rlabel metal2 s 34664 99600 34720 100000 6 io_oeb[27]
port 147 nsew signal output
rlabel metal2 s 35672 99600 35728 100000 6 io_oeb[28]
port 148 nsew signal output
rlabel metal2 s 36680 99600 36736 100000 6 io_oeb[29]
port 149 nsew signal output
rlabel metal2 s 9464 99600 9520 100000 6 io_oeb[2]
port 150 nsew signal output
rlabel metal2 s 37688 99600 37744 100000 6 io_oeb[30]
port 151 nsew signal output
rlabel metal2 s 38696 99600 38752 100000 6 io_oeb[31]
port 152 nsew signal output
rlabel metal2 s 39704 99600 39760 100000 6 io_oeb[32]
port 153 nsew signal output
rlabel metal2 s 40712 99600 40768 100000 6 io_oeb[33]
port 154 nsew signal output
rlabel metal2 s 41720 99600 41776 100000 6 io_oeb[34]
port 155 nsew signal output
rlabel metal2 s 42728 99600 42784 100000 6 io_oeb[35]
port 156 nsew signal output
rlabel metal2 s 43736 99600 43792 100000 6 io_oeb[36]
port 157 nsew signal output
rlabel metal2 s 44744 99600 44800 100000 6 io_oeb[37]
port 158 nsew signal output
rlabel metal2 s 10472 99600 10528 100000 6 io_oeb[3]
port 159 nsew signal output
rlabel metal2 s 11480 99600 11536 100000 6 io_oeb[4]
port 160 nsew signal output
rlabel metal2 s 12488 99600 12544 100000 6 io_oeb[5]
port 161 nsew signal output
rlabel metal2 s 13496 99600 13552 100000 6 io_oeb[6]
port 162 nsew signal output
rlabel metal2 s 14504 99600 14560 100000 6 io_oeb[7]
port 163 nsew signal output
rlabel metal2 s 15512 99600 15568 100000 6 io_oeb[8]
port 164 nsew signal output
rlabel metal2 s 16520 99600 16576 100000 6 io_oeb[9]
port 165 nsew signal output
rlabel metal2 s 7784 99600 7840 100000 6 io_out[0]
port 166 nsew signal output
rlabel metal2 s 17864 99600 17920 100000 6 io_out[10]
port 167 nsew signal output
rlabel metal2 s 18872 99600 18928 100000 6 io_out[11]
port 168 nsew signal output
rlabel metal2 s 19880 99600 19936 100000 6 io_out[12]
port 169 nsew signal output
rlabel metal2 s 20888 99600 20944 100000 6 io_out[13]
port 170 nsew signal output
rlabel metal2 s 21896 99600 21952 100000 6 io_out[14]
port 171 nsew signal output
rlabel metal2 s 22904 99600 22960 100000 6 io_out[15]
port 172 nsew signal output
rlabel metal2 s 23912 99600 23968 100000 6 io_out[16]
port 173 nsew signal output
rlabel metal2 s 24920 99600 24976 100000 6 io_out[17]
port 174 nsew signal output
rlabel metal2 s 25928 99600 25984 100000 6 io_out[18]
port 175 nsew signal output
rlabel metal2 s 26936 99600 26992 100000 6 io_out[19]
port 176 nsew signal output
rlabel metal2 s 8792 99600 8848 100000 6 io_out[1]
port 177 nsew signal output
rlabel metal2 s 27944 99600 28000 100000 6 io_out[20]
port 178 nsew signal output
rlabel metal2 s 28952 99600 29008 100000 6 io_out[21]
port 179 nsew signal output
rlabel metal2 s 29960 99600 30016 100000 6 io_out[22]
port 180 nsew signal output
rlabel metal2 s 30968 99600 31024 100000 6 io_out[23]
port 181 nsew signal output
rlabel metal2 s 31976 99600 32032 100000 6 io_out[24]
port 182 nsew signal output
rlabel metal2 s 32984 99600 33040 100000 6 io_out[25]
port 183 nsew signal output
rlabel metal2 s 33992 99600 34048 100000 6 io_out[26]
port 184 nsew signal output
rlabel metal2 s 35000 99600 35056 100000 6 io_out[27]
port 185 nsew signal output
rlabel metal2 s 36008 99600 36064 100000 6 io_out[28]
port 186 nsew signal output
rlabel metal2 s 37016 99600 37072 100000 6 io_out[29]
port 187 nsew signal output
rlabel metal2 s 9800 99600 9856 100000 6 io_out[2]
port 188 nsew signal output
rlabel metal2 s 38024 99600 38080 100000 6 io_out[30]
port 189 nsew signal output
rlabel metal2 s 39032 99600 39088 100000 6 io_out[31]
port 190 nsew signal output
rlabel metal2 s 40040 99600 40096 100000 6 io_out[32]
port 191 nsew signal output
rlabel metal2 s 41048 99600 41104 100000 6 io_out[33]
port 192 nsew signal output
rlabel metal2 s 42056 99600 42112 100000 6 io_out[34]
port 193 nsew signal output
rlabel metal2 s 43064 99600 43120 100000 6 io_out[35]
port 194 nsew signal output
rlabel metal2 s 44072 99600 44128 100000 6 io_out[36]
port 195 nsew signal output
rlabel metal2 s 45080 99600 45136 100000 6 io_out[37]
port 196 nsew signal output
rlabel metal2 s 10808 99600 10864 100000 6 io_out[3]
port 197 nsew signal output
rlabel metal2 s 11816 99600 11872 100000 6 io_out[4]
port 198 nsew signal output
rlabel metal2 s 12824 99600 12880 100000 6 io_out[5]
port 199 nsew signal output
rlabel metal2 s 13832 99600 13888 100000 6 io_out[6]
port 200 nsew signal output
rlabel metal2 s 14840 99600 14896 100000 6 io_out[7]
port 201 nsew signal output
rlabel metal2 s 15848 99600 15904 100000 6 io_out[8]
port 202 nsew signal output
rlabel metal2 s 16856 99600 16912 100000 6 io_out[9]
port 203 nsew signal output
rlabel metal2 s 95424 0 95480 400 6 irq[0]
port 204 nsew signal output
rlabel metal2 s 96152 0 96208 400 6 irq[1]
port 205 nsew signal output
rlabel metal2 s 96880 0 96936 400 6 irq[2]
port 206 nsew signal output
rlabel metal2 s 2240 0 2296 400 6 la_data_out[0]
port 207 nsew signal output
rlabel metal2 s 75040 0 75096 400 6 la_data_out[100]
port 208 nsew signal output
rlabel metal2 s 75768 0 75824 400 6 la_data_out[101]
port 209 nsew signal output
rlabel metal2 s 76496 0 76552 400 6 la_data_out[102]
port 210 nsew signal output
rlabel metal2 s 77224 0 77280 400 6 la_data_out[103]
port 211 nsew signal output
rlabel metal2 s 77952 0 78008 400 6 la_data_out[104]
port 212 nsew signal output
rlabel metal2 s 78680 0 78736 400 6 la_data_out[105]
port 213 nsew signal output
rlabel metal2 s 79408 0 79464 400 6 la_data_out[106]
port 214 nsew signal output
rlabel metal2 s 80136 0 80192 400 6 la_data_out[107]
port 215 nsew signal output
rlabel metal2 s 80864 0 80920 400 6 la_data_out[108]
port 216 nsew signal output
rlabel metal2 s 81592 0 81648 400 6 la_data_out[109]
port 217 nsew signal output
rlabel metal2 s 9520 0 9576 400 6 la_data_out[10]
port 218 nsew signal output
rlabel metal2 s 82320 0 82376 400 6 la_data_out[110]
port 219 nsew signal output
rlabel metal2 s 83048 0 83104 400 6 la_data_out[111]
port 220 nsew signal output
rlabel metal2 s 83776 0 83832 400 6 la_data_out[112]
port 221 nsew signal output
rlabel metal2 s 84504 0 84560 400 6 la_data_out[113]
port 222 nsew signal output
rlabel metal2 s 85232 0 85288 400 6 la_data_out[114]
port 223 nsew signal output
rlabel metal2 s 85960 0 86016 400 6 la_data_out[115]
port 224 nsew signal output
rlabel metal2 s 86688 0 86744 400 6 la_data_out[116]
port 225 nsew signal output
rlabel metal2 s 87416 0 87472 400 6 la_data_out[117]
port 226 nsew signal output
rlabel metal2 s 88144 0 88200 400 6 la_data_out[118]
port 227 nsew signal output
rlabel metal2 s 88872 0 88928 400 6 la_data_out[119]
port 228 nsew signal output
rlabel metal2 s 10248 0 10304 400 6 la_data_out[11]
port 229 nsew signal output
rlabel metal2 s 89600 0 89656 400 6 la_data_out[120]
port 230 nsew signal output
rlabel metal2 s 90328 0 90384 400 6 la_data_out[121]
port 231 nsew signal output
rlabel metal2 s 91056 0 91112 400 6 la_data_out[122]
port 232 nsew signal output
rlabel metal2 s 91784 0 91840 400 6 la_data_out[123]
port 233 nsew signal output
rlabel metal2 s 92512 0 92568 400 6 la_data_out[124]
port 234 nsew signal output
rlabel metal2 s 93240 0 93296 400 6 la_data_out[125]
port 235 nsew signal output
rlabel metal2 s 93968 0 94024 400 6 la_data_out[126]
port 236 nsew signal output
rlabel metal2 s 94696 0 94752 400 6 la_data_out[127]
port 237 nsew signal output
rlabel metal2 s 10976 0 11032 400 6 la_data_out[12]
port 238 nsew signal output
rlabel metal2 s 11704 0 11760 400 6 la_data_out[13]
port 239 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 la_data_out[14]
port 240 nsew signal output
rlabel metal2 s 13160 0 13216 400 6 la_data_out[15]
port 241 nsew signal output
rlabel metal2 s 13888 0 13944 400 6 la_data_out[16]
port 242 nsew signal output
rlabel metal2 s 14616 0 14672 400 6 la_data_out[17]
port 243 nsew signal output
rlabel metal2 s 15344 0 15400 400 6 la_data_out[18]
port 244 nsew signal output
rlabel metal2 s 16072 0 16128 400 6 la_data_out[19]
port 245 nsew signal output
rlabel metal2 s 2968 0 3024 400 6 la_data_out[1]
port 246 nsew signal output
rlabel metal2 s 16800 0 16856 400 6 la_data_out[20]
port 247 nsew signal output
rlabel metal2 s 17528 0 17584 400 6 la_data_out[21]
port 248 nsew signal output
rlabel metal2 s 18256 0 18312 400 6 la_data_out[22]
port 249 nsew signal output
rlabel metal2 s 18984 0 19040 400 6 la_data_out[23]
port 250 nsew signal output
rlabel metal2 s 19712 0 19768 400 6 la_data_out[24]
port 251 nsew signal output
rlabel metal2 s 20440 0 20496 400 6 la_data_out[25]
port 252 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 la_data_out[26]
port 253 nsew signal output
rlabel metal2 s 21896 0 21952 400 6 la_data_out[27]
port 254 nsew signal output
rlabel metal2 s 22624 0 22680 400 6 la_data_out[28]
port 255 nsew signal output
rlabel metal2 s 23352 0 23408 400 6 la_data_out[29]
port 256 nsew signal output
rlabel metal2 s 3696 0 3752 400 6 la_data_out[2]
port 257 nsew signal output
rlabel metal2 s 24080 0 24136 400 6 la_data_out[30]
port 258 nsew signal output
rlabel metal2 s 24808 0 24864 400 6 la_data_out[31]
port 259 nsew signal output
rlabel metal2 s 25536 0 25592 400 6 la_data_out[32]
port 260 nsew signal output
rlabel metal2 s 26264 0 26320 400 6 la_data_out[33]
port 261 nsew signal output
rlabel metal2 s 26992 0 27048 400 6 la_data_out[34]
port 262 nsew signal output
rlabel metal2 s 27720 0 27776 400 6 la_data_out[35]
port 263 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 la_data_out[36]
port 264 nsew signal output
rlabel metal2 s 29176 0 29232 400 6 la_data_out[37]
port 265 nsew signal output
rlabel metal2 s 29904 0 29960 400 6 la_data_out[38]
port 266 nsew signal output
rlabel metal2 s 30632 0 30688 400 6 la_data_out[39]
port 267 nsew signal output
rlabel metal2 s 4424 0 4480 400 6 la_data_out[3]
port 268 nsew signal output
rlabel metal2 s 31360 0 31416 400 6 la_data_out[40]
port 269 nsew signal output
rlabel metal2 s 32088 0 32144 400 6 la_data_out[41]
port 270 nsew signal output
rlabel metal2 s 32816 0 32872 400 6 la_data_out[42]
port 271 nsew signal output
rlabel metal2 s 33544 0 33600 400 6 la_data_out[43]
port 272 nsew signal output
rlabel metal2 s 34272 0 34328 400 6 la_data_out[44]
port 273 nsew signal output
rlabel metal2 s 35000 0 35056 400 6 la_data_out[45]
port 274 nsew signal output
rlabel metal2 s 35728 0 35784 400 6 la_data_out[46]
port 275 nsew signal output
rlabel metal2 s 36456 0 36512 400 6 la_data_out[47]
port 276 nsew signal output
rlabel metal2 s 37184 0 37240 400 6 la_data_out[48]
port 277 nsew signal output
rlabel metal2 s 37912 0 37968 400 6 la_data_out[49]
port 278 nsew signal output
rlabel metal2 s 5152 0 5208 400 6 la_data_out[4]
port 279 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 la_data_out[50]
port 280 nsew signal output
rlabel metal2 s 39368 0 39424 400 6 la_data_out[51]
port 281 nsew signal output
rlabel metal2 s 40096 0 40152 400 6 la_data_out[52]
port 282 nsew signal output
rlabel metal2 s 40824 0 40880 400 6 la_data_out[53]
port 283 nsew signal output
rlabel metal2 s 41552 0 41608 400 6 la_data_out[54]
port 284 nsew signal output
rlabel metal2 s 42280 0 42336 400 6 la_data_out[55]
port 285 nsew signal output
rlabel metal2 s 43008 0 43064 400 6 la_data_out[56]
port 286 nsew signal output
rlabel metal2 s 43736 0 43792 400 6 la_data_out[57]
port 287 nsew signal output
rlabel metal2 s 44464 0 44520 400 6 la_data_out[58]
port 288 nsew signal output
rlabel metal2 s 45192 0 45248 400 6 la_data_out[59]
port 289 nsew signal output
rlabel metal2 s 5880 0 5936 400 6 la_data_out[5]
port 290 nsew signal output
rlabel metal2 s 45920 0 45976 400 6 la_data_out[60]
port 291 nsew signal output
rlabel metal2 s 46648 0 46704 400 6 la_data_out[61]
port 292 nsew signal output
rlabel metal2 s 47376 0 47432 400 6 la_data_out[62]
port 293 nsew signal output
rlabel metal2 s 48104 0 48160 400 6 la_data_out[63]
port 294 nsew signal output
rlabel metal2 s 48832 0 48888 400 6 la_data_out[64]
port 295 nsew signal output
rlabel metal2 s 49560 0 49616 400 6 la_data_out[65]
port 296 nsew signal output
rlabel metal2 s 50288 0 50344 400 6 la_data_out[66]
port 297 nsew signal output
rlabel metal2 s 51016 0 51072 400 6 la_data_out[67]
port 298 nsew signal output
rlabel metal2 s 51744 0 51800 400 6 la_data_out[68]
port 299 nsew signal output
rlabel metal2 s 52472 0 52528 400 6 la_data_out[69]
port 300 nsew signal output
rlabel metal2 s 6608 0 6664 400 6 la_data_out[6]
port 301 nsew signal output
rlabel metal2 s 53200 0 53256 400 6 la_data_out[70]
port 302 nsew signal output
rlabel metal2 s 53928 0 53984 400 6 la_data_out[71]
port 303 nsew signal output
rlabel metal2 s 54656 0 54712 400 6 la_data_out[72]
port 304 nsew signal output
rlabel metal2 s 55384 0 55440 400 6 la_data_out[73]
port 305 nsew signal output
rlabel metal2 s 56112 0 56168 400 6 la_data_out[74]
port 306 nsew signal output
rlabel metal2 s 56840 0 56896 400 6 la_data_out[75]
port 307 nsew signal output
rlabel metal2 s 57568 0 57624 400 6 la_data_out[76]
port 308 nsew signal output
rlabel metal2 s 58296 0 58352 400 6 la_data_out[77]
port 309 nsew signal output
rlabel metal2 s 59024 0 59080 400 6 la_data_out[78]
port 310 nsew signal output
rlabel metal2 s 59752 0 59808 400 6 la_data_out[79]
port 311 nsew signal output
rlabel metal2 s 7336 0 7392 400 6 la_data_out[7]
port 312 nsew signal output
rlabel metal2 s 60480 0 60536 400 6 la_data_out[80]
port 313 nsew signal output
rlabel metal2 s 61208 0 61264 400 6 la_data_out[81]
port 314 nsew signal output
rlabel metal2 s 61936 0 61992 400 6 la_data_out[82]
port 315 nsew signal output
rlabel metal2 s 62664 0 62720 400 6 la_data_out[83]
port 316 nsew signal output
rlabel metal2 s 63392 0 63448 400 6 la_data_out[84]
port 317 nsew signal output
rlabel metal2 s 64120 0 64176 400 6 la_data_out[85]
port 318 nsew signal output
rlabel metal2 s 64848 0 64904 400 6 la_data_out[86]
port 319 nsew signal output
rlabel metal2 s 65576 0 65632 400 6 la_data_out[87]
port 320 nsew signal output
rlabel metal2 s 66304 0 66360 400 6 la_data_out[88]
port 321 nsew signal output
rlabel metal2 s 67032 0 67088 400 6 la_data_out[89]
port 322 nsew signal output
rlabel metal2 s 8064 0 8120 400 6 la_data_out[8]
port 323 nsew signal output
rlabel metal2 s 67760 0 67816 400 6 la_data_out[90]
port 324 nsew signal output
rlabel metal2 s 68488 0 68544 400 6 la_data_out[91]
port 325 nsew signal output
rlabel metal2 s 69216 0 69272 400 6 la_data_out[92]
port 326 nsew signal output
rlabel metal2 s 69944 0 70000 400 6 la_data_out[93]
port 327 nsew signal output
rlabel metal2 s 70672 0 70728 400 6 la_data_out[94]
port 328 nsew signal output
rlabel metal2 s 71400 0 71456 400 6 la_data_out[95]
port 329 nsew signal output
rlabel metal2 s 72128 0 72184 400 6 la_data_out[96]
port 330 nsew signal output
rlabel metal2 s 72856 0 72912 400 6 la_data_out[97]
port 331 nsew signal output
rlabel metal2 s 73584 0 73640 400 6 la_data_out[98]
port 332 nsew signal output
rlabel metal2 s 74312 0 74368 400 6 la_data_out[99]
port 333 nsew signal output
rlabel metal2 s 8792 0 8848 400 6 la_data_out[9]
port 334 nsew signal output
rlabel metal2 s 99064 0 99120 400 6 reset
port 335 nsew signal output
rlabel metal2 s 98336 0 98392 400 6 start
port 336 nsew signal output
rlabel metal2 s 45752 99600 45808 100000 6 uP_data_mem_addr[0]
port 337 nsew signal input
rlabel metal2 s 47096 99600 47152 100000 6 uP_data_mem_addr[1]
port 338 nsew signal input
rlabel metal2 s 48440 99600 48496 100000 6 uP_data_mem_addr[2]
port 339 nsew signal input
rlabel metal2 s 49784 99600 49840 100000 6 uP_data_mem_addr[3]
port 340 nsew signal input
rlabel metal2 s 51128 99600 51184 100000 6 uP_data_mem_addr[4]
port 341 nsew signal input
rlabel metal2 s 52472 99600 52528 100000 6 uP_data_mem_addr[5]
port 342 nsew signal input
rlabel metal2 s 53816 99600 53872 100000 6 uP_data_mem_addr[6]
port 343 nsew signal input
rlabel metal2 s 55160 99600 55216 100000 6 uP_data_mem_addr[7]
port 344 nsew signal input
rlabel metal2 s 45416 99600 45472 100000 6 uP_dataw_en
port 345 nsew signal input
rlabel metal2 s 46088 99600 46144 100000 6 uP_instr[0]
port 346 nsew signal output
rlabel metal2 s 58520 99600 58576 100000 6 uP_instr[10]
port 347 nsew signal output
rlabel metal2 s 59528 99600 59584 100000 6 uP_instr[11]
port 348 nsew signal output
rlabel metal2 s 60536 99600 60592 100000 6 uP_instr[12]
port 349 nsew signal output
rlabel metal2 s 61544 99600 61600 100000 6 uP_instr[13]
port 350 nsew signal output
rlabel metal2 s 62216 99600 62272 100000 6 uP_instr[14]
port 351 nsew signal output
rlabel metal2 s 62888 99600 62944 100000 6 uP_instr[15]
port 352 nsew signal output
rlabel metal2 s 47432 99600 47488 100000 6 uP_instr[1]
port 353 nsew signal output
rlabel metal2 s 48776 99600 48832 100000 6 uP_instr[2]
port 354 nsew signal output
rlabel metal2 s 50120 99600 50176 100000 6 uP_instr[3]
port 355 nsew signal output
rlabel metal2 s 51464 99600 51520 100000 6 uP_instr[4]
port 356 nsew signal output
rlabel metal2 s 52808 99600 52864 100000 6 uP_instr[5]
port 357 nsew signal output
rlabel metal2 s 54152 99600 54208 100000 6 uP_instr[6]
port 358 nsew signal output
rlabel metal2 s 55496 99600 55552 100000 6 uP_instr[7]
port 359 nsew signal output
rlabel metal2 s 56504 99600 56560 100000 6 uP_instr[8]
port 360 nsew signal output
rlabel metal2 s 57512 99600 57568 100000 6 uP_instr[9]
port 361 nsew signal output
rlabel metal2 s 46424 99600 46480 100000 6 uP_instr_mem_addr[0]
port 362 nsew signal input
rlabel metal2 s 58856 99600 58912 100000 6 uP_instr_mem_addr[10]
port 363 nsew signal input
rlabel metal2 s 59864 99600 59920 100000 6 uP_instr_mem_addr[11]
port 364 nsew signal input
rlabel metal2 s 60872 99600 60928 100000 6 uP_instr_mem_addr[12]
port 365 nsew signal input
rlabel metal2 s 47768 99600 47824 100000 6 uP_instr_mem_addr[1]
port 366 nsew signal input
rlabel metal2 s 49112 99600 49168 100000 6 uP_instr_mem_addr[2]
port 367 nsew signal input
rlabel metal2 s 50456 99600 50512 100000 6 uP_instr_mem_addr[3]
port 368 nsew signal input
rlabel metal2 s 51800 99600 51856 100000 6 uP_instr_mem_addr[4]
port 369 nsew signal input
rlabel metal2 s 53144 99600 53200 100000 6 uP_instr_mem_addr[5]
port 370 nsew signal input
rlabel metal2 s 54488 99600 54544 100000 6 uP_instr_mem_addr[6]
port 371 nsew signal input
rlabel metal2 s 55832 99600 55888 100000 6 uP_instr_mem_addr[7]
port 372 nsew signal input
rlabel metal2 s 56840 99600 56896 100000 6 uP_instr_mem_addr[8]
port 373 nsew signal input
rlabel metal2 s 57848 99600 57904 100000 6 uP_instr_mem_addr[9]
port 374 nsew signal input
rlabel metal2 s 46760 99600 46816 100000 6 uP_write_data[0]
port 375 nsew signal input
rlabel metal2 s 59192 99600 59248 100000 6 uP_write_data[10]
port 376 nsew signal input
rlabel metal2 s 60200 99600 60256 100000 6 uP_write_data[11]
port 377 nsew signal input
rlabel metal2 s 61208 99600 61264 100000 6 uP_write_data[12]
port 378 nsew signal input
rlabel metal2 s 61880 99600 61936 100000 6 uP_write_data[13]
port 379 nsew signal input
rlabel metal2 s 62552 99600 62608 100000 6 uP_write_data[14]
port 380 nsew signal input
rlabel metal2 s 63224 99600 63280 100000 6 uP_write_data[15]
port 381 nsew signal input
rlabel metal2 s 48104 99600 48160 100000 6 uP_write_data[1]
port 382 nsew signal input
rlabel metal2 s 49448 99600 49504 100000 6 uP_write_data[2]
port 383 nsew signal input
rlabel metal2 s 50792 99600 50848 100000 6 uP_write_data[3]
port 384 nsew signal input
rlabel metal2 s 52136 99600 52192 100000 6 uP_write_data[4]
port 385 nsew signal input
rlabel metal2 s 53480 99600 53536 100000 6 uP_write_data[5]
port 386 nsew signal input
rlabel metal2 s 54824 99600 54880 100000 6 uP_write_data[6]
port 387 nsew signal input
rlabel metal2 s 56168 99600 56224 100000 6 uP_write_data[7]
port 388 nsew signal input
rlabel metal2 s 57176 99600 57232 100000 6 uP_write_data[8]
port 389 nsew signal input
rlabel metal2 s 58184 99600 58240 100000 6 uP_write_data[9]
port 390 nsew signal input
rlabel metal4 s 2224 1538 2384 98422 6 vdd
port 391 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 vdd
port 391 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 vdd
port 391 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 vdd
port 391 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 vdd
port 391 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 vdd
port 391 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 98422 6 vdd
port 391 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 vss
port 392 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 vss
port 392 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 vss
port 392 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 vss
port 392 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 vss
port 392 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 vss
port 392 nsew ground bidirectional
rlabel metal2 s 784 0 840 400 6 wb_clk_i
port 393 nsew signal input
rlabel metal2 s 1512 0 1568 400 6 wb_rst_i
port 394 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4985672
string GDS_FILE /home/radhe/tapeout_projects/radhe_gf180nm/openlane/io_interface/runs/22_12_08_14_26/results/signoff/io_interface.magic.gds
string GDS_START 162452
<< end >>

