// This is the unpowered netlist.
module io_interface (Serial_input,
    Serial_output,
    clk,
    data_mem_sel,
    dataw_en,
    hlt,
    instr_mem_sel,
    instrw_en,
    reset,
    start,
    uP_dataw_en,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    data_mem_addr,
    data_read_data,
    data_write_data,
    dataw_en_8bit,
    instr,
    instr_mem_addr,
    instr_write_data,
    instrw_en_8bit,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    uP_data_mem_addr,
    uP_instr,
    uP_instr_mem_addr,
    uP_write_data,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input Serial_input;
 output Serial_output;
 output clk;
 output data_mem_sel;
 output dataw_en;
 input hlt;
 output instr_mem_sel;
 output instrw_en;
 output reset;
 output start;
 input uP_dataw_en;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 output [7:0] data_mem_addr;
 input [15:0] data_read_data;
 output [15:0] data_write_data;
 output [7:0] dataw_en_8bit;
 input [15:0] instr;
 output [7:0] instr_mem_addr;
 output [15:0] instr_write_data;
 output [7:0] instrw_en_8bit;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [7:0] uP_data_mem_addr;
 output [15:0] uP_instr;
 input [12:0] uP_instr_mem_addr;
 input [15:0] uP_write_data;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire net713;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire \data_load_addr[0] ;
 wire \data_load_addr[1] ;
 wire \data_load_addr[2] ;
 wire \data_load_addr[3] ;
 wire \data_load_addr[4] ;
 wire \data_load_addr[5] ;
 wire \data_load_addr[6] ;
 wire \data_load_addr[7] ;
 wire net714;
 wire \instr_load_addr[0] ;
 wire \instr_load_addr[10] ;
 wire \instr_load_addr[11] ;
 wire \instr_load_addr[12] ;
 wire \instr_load_addr[1] ;
 wire \instr_load_addr[2] ;
 wire \instr_load_addr[3] ;
 wire \instr_load_addr[4] ;
 wire \instr_load_addr[5] ;
 wire \instr_load_addr[6] ;
 wire \instr_load_addr[7] ;
 wire \instr_load_addr[8] ;
 wire \instr_load_addr[9] ;
 wire net715;
 wire net716;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net717;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net718;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net732;
 wire net778;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0440_ (.I(net34),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0441_ (.I(net51),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0442_ (.I(_0165_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0443_ (.I(net52),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0444_ (.I(_0167_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0445_ (.I0(net1),
    .I1(net18),
    .I2(\data_load_addr[0] ),
    .I3(\instr_load_addr[0] ),
    .S0(_0166_),
    .S1(_0168_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0446_ (.I(net50),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0447_ (.I(_0170_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0448_ (.I0(_0164_),
    .I1(_0169_),
    .S(_0171_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0449_ (.I(_0172_),
    .Z(net482));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0450_ (.I(net35),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0451_ (.I0(net8),
    .I1(net25),
    .I2(\data_load_addr[1] ),
    .I3(\instr_load_addr[1] ),
    .S0(_0166_),
    .S1(_0168_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0452_ (.I0(_0173_),
    .I1(_0174_),
    .S(_0171_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0453_ (.I(_0175_),
    .Z(net489));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0454_ (.I(net36),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0455_ (.I(\data_load_addr[2] ),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0456_ (.I(\instr_load_addr[2] ),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0457_ (.I(net52),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0458_ (.I0(net9),
    .I1(net26),
    .I2(_0177_),
    .I3(_0178_),
    .S0(_0166_),
    .S1(_0179_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0459_ (.I0(_0176_),
    .I1(_0180_),
    .S(_0171_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0460_ (.I(_0181_),
    .Z(net490));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0461_ (.I(net37),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0462_ (.I(_0165_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0463_ (.I0(net10),
    .I1(net27),
    .I2(\data_load_addr[3] ),
    .I3(\instr_load_addr[3] ),
    .S0(_0183_),
    .S1(_0179_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0464_ (.I0(_0182_),
    .I1(_0184_),
    .S(_0171_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0465_ (.I(_0185_),
    .Z(net492));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0466_ (.I(net38),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0467_ (.I(\instr_load_addr[4] ),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0468_ (.I0(net11),
    .I1(net28),
    .I2(\data_load_addr[4] ),
    .I3(_0187_),
    .S0(_0183_),
    .S1(_0179_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0469_ (.I(_0170_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0470_ (.I0(_0186_),
    .I1(_0188_),
    .S(_0189_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0471_ (.I(_0190_),
    .Z(net493));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0472_ (.I(net39),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0473_ (.I0(net12),
    .I1(net29),
    .I2(\data_load_addr[5] ),
    .I3(\instr_load_addr[5] ),
    .S0(_0183_),
    .S1(_0179_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0474_ (.I0(_0191_),
    .I1(_0192_),
    .S(_0189_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0475_ (.I(_0193_),
    .Z(net494));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0476_ (.I(net40),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0477_ (.I(\instr_load_addr[6] ),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0478_ (.I0(net13),
    .I1(net30),
    .I2(\data_load_addr[6] ),
    .I3(_0195_),
    .S0(_0183_),
    .S1(_0167_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0479_ (.I0(_0194_),
    .I1(_0196_),
    .S(_0189_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0480_ (.I(_0197_),
    .Z(net495));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0481_ (.I(net41),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0482_ (.I0(net14),
    .I1(net31),
    .I2(\data_load_addr[7] ),
    .I3(\instr_load_addr[7] ),
    .S0(_0165_),
    .S1(_0167_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0483_ (.I0(_0198_),
    .I1(_0199_),
    .S(_0189_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0484_ (.I(_0200_),
    .Z(net496));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0485_ (.I(net50),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0486_ (.I(_0201_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0487_ (.A1(_0165_),
    .A2(_0167_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0488_ (.I(_0203_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0489_ (.A1(net51),
    .A2(net52),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0490_ (.I(_0205_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0491_ (.I(net51),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0492_ (.A1(_0207_),
    .A2(net52),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0493_ (.I(_0208_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0494_ (.A1(\instr_load_addr[8] ),
    .A2(_0204_),
    .B1(_0206_),
    .B2(net15),
    .C1(_0209_),
    .C2(net32),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0495_ (.I(net50),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0496_ (.A1(_0211_),
    .A2(net699),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0497_ (.A1(_0202_),
    .A2(_0210_),
    .B(_0212_),
    .ZN(net497));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0498_ (.A1(\instr_load_addr[9] ),
    .A2(_0204_),
    .B1(_0206_),
    .B2(net16),
    .C1(_0209_),
    .C2(net33),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0499_ (.A1(_0211_),
    .A2(net698),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0500_ (.A1(_0202_),
    .A2(_0213_),
    .B(_0214_),
    .ZN(net498));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0501_ (.A1(\instr_load_addr[10] ),
    .A2(_0204_),
    .B1(_0206_),
    .B2(net2),
    .C1(_0209_),
    .C2(net19),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0502_ (.A1(_0211_),
    .A2(net697),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0503_ (.A1(_0202_),
    .A2(_0215_),
    .B(_0216_),
    .ZN(net483));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0504_ (.I(_0201_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0505_ (.A1(\instr_load_addr[11] ),
    .A2(_0204_),
    .B1(_0206_),
    .B2(net3),
    .C1(_0209_),
    .C2(net20),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0506_ (.I(_0201_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0507_ (.A1(_0219_),
    .A2(net696),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0508_ (.A1(_0217_),
    .A2(_0218_),
    .B(_0220_),
    .ZN(net484));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0509_ (.A1(\instr_load_addr[12] ),
    .A2(_0203_),
    .B1(_0205_),
    .B2(net4),
    .C1(_0208_),
    .C2(net21),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0510_ (.A1(_0219_),
    .A2(net695),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0511_ (.A1(_0217_),
    .A2(_0221_),
    .B(_0222_),
    .ZN(net485));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0512_ (.I(_0205_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0513_ (.I(_0208_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0514_ (.A1(net5),
    .A2(_0223_),
    .B1(_0224_),
    .B2(net22),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0515_ (.A1(_0219_),
    .A2(net47),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0516_ (.A1(_0217_),
    .A2(_0225_),
    .B(_0226_),
    .ZN(net486));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0517_ (.A1(net6),
    .A2(_0223_),
    .B1(_0224_),
    .B2(net23),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0518_ (.A1(_0219_),
    .A2(net48),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0519_ (.A1(_0217_),
    .A2(_0227_),
    .B(_0228_),
    .ZN(net487));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0520_ (.A1(net7),
    .A2(_0223_),
    .B1(_0224_),
    .B2(net24),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0521_ (.A1(_0201_),
    .A2(net49),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0522_ (.A1(_0211_),
    .A2(_0229_),
    .B(_0230_),
    .ZN(net488));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0523_ (.I(\data_load_addr[0] ),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0524_ (.I(net694),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0525_ (.I(_0232_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0526_ (.I0(_0231_),
    .I1(net309),
    .S(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0527_ (.I(_0234_),
    .Z(net416));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0528_ (.I(\data_load_addr[1] ),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0529_ (.I0(_0235_),
    .I1(net310),
    .S(_0233_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0530_ (.I(_0236_),
    .Z(net417));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0531_ (.I(net694),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0532_ (.I(_0237_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0533_ (.I0(_0177_),
    .I1(net311),
    .S(_0238_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0534_ (.I(_0239_),
    .Z(net418));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0535_ (.I0(\data_load_addr[3] ),
    .I1(net312),
    .S(_0238_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0536_ (.I(_0240_),
    .Z(net419));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0537_ (.I0(\data_load_addr[4] ),
    .I1(net313),
    .S(_0238_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0538_ (.I(_0241_),
    .Z(net420));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0539_ (.I(\data_load_addr[5] ),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0540_ (.I0(_0242_),
    .I1(net314),
    .S(_0238_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0541_ (.I(_0243_),
    .Z(net421));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0542_ (.I(net694),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0543_ (.I(_0244_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0544_ (.I0(\data_load_addr[6] ),
    .I1(net315),
    .S(_0245_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0545_ (.I(_0246_),
    .Z(net422));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0546_ (.I0(\data_load_addr[7] ),
    .I1(net316),
    .S(_0245_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0547_ (.I(_0247_),
    .Z(net423));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0548_ (.I(\instr_load_addr[0] ),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0549_ (.I0(_0248_),
    .I1(net318),
    .S(_0245_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0550_ (.I(_0249_),
    .Z(net449));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0551_ (.I(\instr_load_addr[1] ),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0552_ (.I0(_0250_),
    .I1(net319),
    .S(_0245_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0553_ (.I(_0251_),
    .Z(net450));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0554_ (.I(_0244_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0555_ (.I0(_0178_),
    .I1(net320),
    .S(_0252_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0556_ (.I(_0253_),
    .Z(net451));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0557_ (.I0(\instr_load_addr[3] ),
    .I1(net321),
    .S(_0252_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0558_ (.I(_0254_),
    .Z(net452));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0559_ (.I0(_0187_),
    .I1(net322),
    .S(_0252_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0560_ (.I(_0255_),
    .Z(net453));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0561_ (.I0(\instr_load_addr[5] ),
    .I1(net323),
    .S(_0252_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0562_ (.I(_0256_),
    .Z(net454));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0563_ (.I(_0244_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0564_ (.I0(_0195_),
    .I1(net324),
    .S(_0257_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0565_ (.I(_0258_),
    .Z(net455));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0566_ (.I0(\instr_load_addr[7] ),
    .I1(net325),
    .S(_0257_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0567_ (.I(_0259_),
    .Z(net456));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0568_ (.I(_0237_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0569_ (.A1(net18),
    .A2(_0260_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0570_ (.I(_0261_),
    .Z(net627));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0571_ (.A1(net25),
    .A2(_0260_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0572_ (.I(_0262_),
    .Z(net634));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0573_ (.I(net26),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0574_ (.I(_0232_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0575_ (.I(_0264_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0576_ (.A1(_0263_),
    .A2(_0265_),
    .ZN(net635));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0577_ (.A1(net27),
    .A2(_0260_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0578_ (.I(_0266_),
    .Z(net636));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0579_ (.A1(net28),
    .A2(_0260_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0580_ (.I(_0267_),
    .Z(net637));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0581_ (.I(_0237_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0582_ (.A1(net29),
    .A2(_0268_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0583_ (.I(_0269_),
    .Z(net638));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0584_ (.A1(net30),
    .A2(_0268_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0585_ (.I(_0270_),
    .Z(net639));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0586_ (.A1(net31),
    .A2(_0268_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0587_ (.I(_0271_),
    .Z(net640));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0588_ (.A1(net32),
    .A2(_0268_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0589_ (.I(_0272_),
    .Z(net641));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0590_ (.I(_0237_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0591_ (.A1(net33),
    .A2(_0273_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0592_ (.I(_0274_),
    .Z(net642));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0593_ (.A1(net19),
    .A2(_0273_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0594_ (.I(_0275_),
    .Z(net628));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0595_ (.A1(net20),
    .A2(_0273_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0596_ (.I(_0276_),
    .Z(net629));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0597_ (.A1(net21),
    .A2(_0273_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0598_ (.I(_0277_),
    .Z(net630));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0599_ (.I(net22),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0600_ (.A1(_0278_),
    .A2(_0265_),
    .ZN(net631));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0601_ (.A1(net23),
    .A2(_0233_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0602_ (.I(_0279_),
    .Z(net632));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0603_ (.A1(net24),
    .A2(_0233_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0604_ (.I(_0280_),
    .Z(net633));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0605_ (.A1(_0170_),
    .A2(net694),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0606_ (.A1(_0265_),
    .A2(net317),
    .B1(_0223_),
    .B2(_0281_),
    .ZN(net440));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0607_ (.I0(net34),
    .I1(net326),
    .S(_0257_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0608_ (.I(_0282_),
    .Z(net424));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0609_ (.I0(net35),
    .I1(net333),
    .S(_0257_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0610_ (.I(_0283_),
    .Z(net431));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0611_ (.I(_0244_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0612_ (.I0(net36),
    .I1(net334),
    .S(_0284_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0613_ (.I(_0285_),
    .Z(net432));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0614_ (.I0(net37),
    .I1(net335),
    .S(_0284_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0615_ (.I(_0286_),
    .Z(net433));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0616_ (.I0(net38),
    .I1(net336),
    .S(_0284_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0617_ (.I(_0287_),
    .Z(net434));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0618_ (.I0(net39),
    .I1(net337),
    .S(_0284_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0619_ (.I(_0288_),
    .Z(net435));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0620_ (.I(_0232_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0621_ (.I0(net40),
    .I1(net338),
    .S(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0622_ (.I(_0290_),
    .Z(net436));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0623_ (.I0(net41),
    .I1(net339),
    .S(_0289_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0624_ (.I(_0291_),
    .Z(net437));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0625_ (.I0(net699),
    .I1(net340),
    .S(_0289_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0626_ (.I(_0292_),
    .Z(net438));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0627_ (.I0(net698),
    .I1(net341),
    .S(_0289_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0628_ (.I(_0293_),
    .Z(net439));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0629_ (.I(_0232_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0630_ (.I0(net697),
    .I1(net327),
    .S(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0631_ (.I(_0295_),
    .Z(net425));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0632_ (.I0(net696),
    .I1(net328),
    .S(_0294_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0633_ (.I(_0296_),
    .Z(net426));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0634_ (.I0(net695),
    .I1(net329),
    .S(_0294_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0635_ (.I(_0297_),
    .Z(net427));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0636_ (.I0(net47),
    .I1(net330),
    .S(_0294_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0637_ (.I(_0298_),
    .Z(net428));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0638_ (.I0(net48),
    .I1(net331),
    .S(_0264_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0639_ (.I(_0299_),
    .Z(net429));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0640_ (.I0(net49),
    .I1(net332),
    .S(_0264_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0641_ (.I(_0300_),
    .Z(net430));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0642_ (.A1(net292),
    .A2(net291),
    .A3(net294),
    .A4(net293),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0643_ (.A1(net288),
    .A2(net287),
    .A3(net290),
    .A4(net289),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0644_ (.A1(net296),
    .A2(net295),
    .A3(net299),
    .A4(net298),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0645_ (.A1(net301),
    .A2(net300),
    .A3(net303),
    .A4(net302),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0646_ (.A1(_0301_),
    .A2(_0302_),
    .A3(_0303_),
    .A4(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0647_ (.A1(net274),
    .A2(net273),
    .A3(net277),
    .A4(net276),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0648_ (.A1(net270),
    .A2(net269),
    .A3(net272),
    .A4(net271),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0649_ (.A1(net279),
    .A2(net278),
    .A3(net281),
    .A4(net280),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0650_ (.A1(net283),
    .A2(net282),
    .A3(net285),
    .A4(net284),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0651_ (.A1(_0306_),
    .A2(_0307_),
    .A3(_0308_),
    .A4(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0652_ (.A1(net183),
    .A2(net182),
    .A3(net185),
    .A4(net184),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0653_ (.A1(net305),
    .A2(net304),
    .A3(net307),
    .A4(net306),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0654_ (.A1(net187),
    .A2(net186),
    .A3(net189),
    .A4(net188),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0655_ (.A1(net191),
    .A2(net190),
    .A3(net194),
    .A4(net193),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0656_ (.A1(_0311_),
    .A2(_0312_),
    .A3(_0313_),
    .A4(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0657_ (.A1(net200),
    .A2(net199),
    .A3(net202),
    .A4(net201),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0658_ (.A1(net196),
    .A2(net195),
    .A3(net198),
    .A4(net197),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0659_ (.A1(net205),
    .A2(net204),
    .A3(net207),
    .A4(net206),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0660_ (.A1(net209),
    .A2(net208),
    .A3(net211),
    .A4(net210),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0661_ (.A1(_0316_),
    .A2(_0317_),
    .A3(_0318_),
    .A4(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0662_ (.A1(_0305_),
    .A2(_0310_),
    .A3(_0315_),
    .A4(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0663_ (.A1(net222),
    .A2(net221),
    .A3(net224),
    .A4(net223),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0664_ (.A1(net217),
    .A2(net216),
    .A3(net219),
    .A4(net218),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0665_ (.A1(net226),
    .A2(net225),
    .A3(net228),
    .A4(net227),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0666_ (.A1(net230),
    .A2(net229),
    .A3(net233),
    .A4(net232),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0667_ (.A1(_0322_),
    .A2(_0323_),
    .A3(_0324_),
    .A4(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0668_ (.A1(net242),
    .A2(net231),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0669_ (.A1(net264),
    .A2(net253),
    .A3(net286),
    .A4(net275),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0670_ (.A1(net213),
    .A2(net212),
    .A3(net215),
    .A4(net214),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0671_ (.A1(net308),
    .A2(net297),
    .A3(net203),
    .A4(net192),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0672_ (.A1(_0327_),
    .A2(_0328_),
    .A3(_0329_),
    .A4(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0673_ (.A1(net257),
    .A2(net256),
    .A3(net259),
    .A4(net258),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0674_ (.A1(net252),
    .A2(net251),
    .A3(net255),
    .A4(net254),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0675_ (.A1(net261),
    .A2(net260),
    .A3(net263),
    .A4(net262),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0676_ (.A1(net266),
    .A2(net265),
    .A3(net268),
    .A4(net267),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0677_ (.A1(_0332_),
    .A2(_0333_),
    .A3(_0334_),
    .A4(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0678_ (.A1(net239),
    .A2(net238),
    .A3(net241),
    .A4(net240),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0679_ (.A1(net235),
    .A2(net234),
    .A3(net237),
    .A4(net236),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0680_ (.A1(net244),
    .A2(net243),
    .A3(net246),
    .A4(net245),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0681_ (.A1(net248),
    .A2(net247),
    .A3(net250),
    .A4(net249),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0682_ (.A1(_0337_),
    .A2(_0338_),
    .A3(_0339_),
    .A4(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0683_ (.A1(_0326_),
    .A2(_0331_),
    .A3(_0336_),
    .A4(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0684_ (.A1(_0321_),
    .A2(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0685_ (.I(_0343_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0686_ (.I(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0687_ (.A1(net104),
    .A2(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0688_ (.I(_0346_),
    .Z(net547));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0689_ (.I(_0343_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0690_ (.I(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0691_ (.I0(net409),
    .I1(net115),
    .S(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0692_ (.I(_0349_),
    .Z(net558));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0693_ (.I0(net410),
    .I1(net126),
    .S(_0348_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0694_ (.I(_0350_),
    .Z(net569));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0695_ (.I0(net411),
    .I1(net137),
    .S(_0348_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0696_ (.I(_0351_),
    .Z(net580));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0697_ (.I(_0347_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0698_ (.I(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0699_ (.I0(net412),
    .I1(net148),
    .S(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0700_ (.I(_0354_),
    .Z(net591));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0701_ (.I0(net414),
    .I1(net159),
    .S(_0353_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0702_ (.I(_0355_),
    .Z(net602));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0703_ (.I0(net376),
    .I1(net170),
    .S(_0353_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0704_ (.I(_0356_),
    .Z(net613));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0705_ (.I0(net413),
    .I1(net181),
    .S(_0353_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0706_ (.I(_0357_),
    .Z(net624));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0707_ (.I(_0352_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0708_ (.I0(net365),
    .I1(net65),
    .S(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0709_ (.I(_0359_),
    .Z(net509));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0710_ (.I0(net367),
    .I1(net76),
    .S(_0358_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0711_ (.I(_0360_),
    .Z(net520));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0712_ (.I0(net368),
    .I1(net85),
    .S(_0358_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0713_ (.I(_0361_),
    .Z(net529));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0714_ (.A1(net86),
    .A2(_0345_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0715_ (.I(_0362_),
    .Z(net530));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0716_ (.A1(net87),
    .A2(_0345_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0717_ (.I(_0363_),
    .Z(net531));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0718_ (.A1(net88),
    .A2(_0345_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0719_ (.I(_0364_),
    .Z(net532));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0720_ (.I0(net627),
    .I1(net89),
    .S(_0358_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0721_ (.I(_0365_),
    .Z(net533));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0722_ (.I(_0352_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0723_ (.I0(net634),
    .I1(net90),
    .S(_0366_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0724_ (.I(_0367_),
    .Z(net534));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0725_ (.I0(net635),
    .I1(net91),
    .S(_0366_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0726_ (.I(_0368_),
    .Z(net535));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0727_ (.I0(net636),
    .I1(net92),
    .S(_0366_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0728_ (.I(_0369_),
    .Z(net536));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0729_ (.I0(net637),
    .I1(net94),
    .S(_0366_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0730_ (.I(_0370_),
    .Z(net537));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0731_ (.I(_0352_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0732_ (.I0(net638),
    .I1(net95),
    .S(_0371_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0733_ (.I(_0372_),
    .Z(net538));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0734_ (.I0(net639),
    .I1(net96),
    .S(_0371_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0735_ (.I(_0373_),
    .Z(net539));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0736_ (.I0(net640),
    .I1(net97),
    .S(_0371_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0737_ (.I(_0374_),
    .Z(net540));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0738_ (.I0(net641),
    .I1(net98),
    .S(_0371_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0739_ (.I(_0375_),
    .Z(net541));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0740_ (.I(_0347_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0741_ (.I(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0742_ (.I0(net642),
    .I1(net99),
    .S(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0743_ (.I(_0378_),
    .Z(net542));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0744_ (.I0(net628),
    .I1(net100),
    .S(_0377_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0745_ (.I(_0379_),
    .Z(net543));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0746_ (.I0(net629),
    .I1(net101),
    .S(_0377_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0747_ (.I(_0380_),
    .Z(net544));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0748_ (.I0(net630),
    .I1(net102),
    .S(_0377_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0749_ (.I(_0381_),
    .Z(net545));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0750_ (.I(_0376_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0751_ (.I0(net631),
    .I1(net103),
    .S(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0752_ (.I(_0383_),
    .Z(net546));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0753_ (.I0(net632),
    .I1(net105),
    .S(_0382_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0754_ (.I(_0384_),
    .Z(net548));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0755_ (.I0(net633),
    .I1(net106),
    .S(_0382_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0756_ (.I(_0385_),
    .Z(net549));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0757_ (.I0(net449),
    .I1(net107),
    .S(_0382_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0758_ (.I(_0386_),
    .Z(net550));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0759_ (.I(_0376_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0760_ (.I0(net450),
    .I1(net108),
    .S(_0387_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0761_ (.I(_0388_),
    .Z(net551));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0762_ (.I0(net451),
    .I1(net109),
    .S(_0387_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0763_ (.I(_0389_),
    .Z(net552));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0764_ (.I0(net452),
    .I1(net110),
    .S(_0387_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0765_ (.I(_0390_),
    .Z(net553));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0766_ (.I0(net453),
    .I1(net111),
    .S(_0387_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0767_ (.I(_0391_),
    .Z(net554));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0768_ (.I(_0376_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0769_ (.I0(net454),
    .I1(net112),
    .S(_0392_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0770_ (.I(_0393_),
    .Z(net555));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0771_ (.I0(net455),
    .I1(net113),
    .S(_0392_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0772_ (.I(_0394_),
    .Z(net556));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0773_ (.I0(net456),
    .I1(net114),
    .S(_0392_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0774_ (.I(_0395_),
    .Z(net557));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0775_ (.I(_0344_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0776_ (.A1(net116),
    .A2(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0777_ (.I(_0397_),
    .Z(net559));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0778_ (.A1(net117),
    .A2(_0396_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0779_ (.I(_0398_),
    .Z(net560));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0780_ (.A1(net118),
    .A2(_0396_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0781_ (.I(_0399_),
    .Z(net561));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0782_ (.A1(net119),
    .A2(_0396_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0783_ (.I(_0400_),
    .Z(net562));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0784_ (.A1(net120),
    .A2(_0348_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0785_ (.I(_0401_),
    .Z(net563));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0786_ (.I0(net424),
    .I1(net121),
    .S(_0392_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0787_ (.I(_0402_),
    .Z(net564));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0788_ (.I(_0347_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0789_ (.I(_0403_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0790_ (.I0(net431),
    .I1(net122),
    .S(_0404_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0791_ (.I(_0405_),
    .Z(net565));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0792_ (.I0(net432),
    .I1(net123),
    .S(_0404_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0793_ (.I(_0406_),
    .Z(net566));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0794_ (.I0(net433),
    .I1(net124),
    .S(_0404_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0795_ (.I(_0407_),
    .Z(net567));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0796_ (.I0(net434),
    .I1(net125),
    .S(_0404_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0797_ (.I(_0408_),
    .Z(net568));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0798_ (.I(_0403_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0799_ (.I0(net435),
    .I1(net127),
    .S(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0800_ (.I(_0410_),
    .Z(net570));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0801_ (.I0(net436),
    .I1(net128),
    .S(_0409_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0802_ (.I(_0411_),
    .Z(net571));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0803_ (.I0(net437),
    .I1(net129),
    .S(_0409_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0804_ (.I(_0412_),
    .Z(net572));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0805_ (.I0(net438),
    .I1(net130),
    .S(_0409_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0806_ (.I(_0413_),
    .Z(net573));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0807_ (.I(_0403_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0808_ (.I0(net439),
    .I1(net131),
    .S(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0809_ (.I(_0415_),
    .Z(net574));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0810_ (.I0(net425),
    .I1(net132),
    .S(_0414_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0811_ (.I(_0416_),
    .Z(net575));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0812_ (.I0(net426),
    .I1(net133),
    .S(_0414_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0813_ (.I(_0417_),
    .Z(net576));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0814_ (.I0(net427),
    .I1(net134),
    .S(_0414_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0815_ (.I(_0418_),
    .Z(net577));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0816_ (.I(_0403_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0817_ (.I0(net428),
    .I1(net135),
    .S(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0818_ (.I(_0420_),
    .Z(net578));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0819_ (.I0(net429),
    .I1(net136),
    .S(_0419_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0820_ (.I(_0421_),
    .Z(net579));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0821_ (.I0(net430),
    .I1(net138),
    .S(_0419_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0822_ (.I(_0422_),
    .Z(net581));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0823_ (.I0(net1),
    .I1(net139),
    .S(_0419_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0824_ (.I(_0423_),
    .Z(net582));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0825_ (.I(_0343_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0826_ (.I(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0827_ (.I(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0828_ (.I0(net8),
    .I1(net140),
    .S(_0426_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0829_ (.I(_0427_),
    .Z(net583));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0830_ (.I0(net9),
    .I1(net141),
    .S(_0426_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0831_ (.I(_0428_),
    .Z(net584));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0832_ (.I0(net10),
    .I1(net142),
    .S(_0426_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0833_ (.I(_0429_),
    .Z(net585));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0834_ (.I0(net11),
    .I1(net143),
    .S(_0426_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0835_ (.I(_0430_),
    .Z(net586));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0836_ (.I(_0425_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0837_ (.I0(net12),
    .I1(net144),
    .S(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0838_ (.I(_0432_),
    .Z(net587));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0839_ (.I0(net13),
    .I1(net145),
    .S(_0431_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0840_ (.I(_0433_),
    .Z(net588));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0841_ (.I0(net14),
    .I1(net146),
    .S(_0431_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0842_ (.I(_0434_),
    .Z(net589));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0843_ (.I0(net15),
    .I1(net147),
    .S(_0431_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0844_ (.I(_0435_),
    .Z(net590));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0845_ (.I(_0425_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0846_ (.I0(net16),
    .I1(net149),
    .S(_0436_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0847_ (.I(_0437_),
    .Z(net592));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0848_ (.I0(net2),
    .I1(net150),
    .S(_0436_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0849_ (.I(_0438_),
    .Z(net593));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0850_ (.I0(net3),
    .I1(net151),
    .S(_0436_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0851_ (.I(_0439_),
    .Z(net594));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0852_ (.I0(net4),
    .I1(net152),
    .S(_0436_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0853_ (.I(_0021_),
    .Z(net595));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0854_ (.I(_0425_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0855_ (.I0(net5),
    .I1(net153),
    .S(_0022_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0856_ (.I(_0023_),
    .Z(net596));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0857_ (.I0(net6),
    .I1(net154),
    .S(_0022_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0858_ (.I(_0024_),
    .Z(net597));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0859_ (.I0(net7),
    .I1(net155),
    .S(_0022_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0860_ (.I(_0025_),
    .Z(net598));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0861_ (.I0(net416),
    .I1(net156),
    .S(_0022_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0862_ (.I(_0026_),
    .Z(net599));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0863_ (.I(_0424_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0864_ (.I(_0027_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0865_ (.I0(net417),
    .I1(net157),
    .S(_0028_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0866_ (.I(_0029_),
    .Z(net600));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0867_ (.I0(net418),
    .I1(net158),
    .S(_0028_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0868_ (.I(_0030_),
    .Z(net601));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0869_ (.I0(net419),
    .I1(net160),
    .S(_0028_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0870_ (.I(_0031_),
    .Z(net603));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0871_ (.I0(net420),
    .I1(net161),
    .S(_0028_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0872_ (.I(_0032_),
    .Z(net604));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0873_ (.I(_0027_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0874_ (.I0(net421),
    .I1(net162),
    .S(_0033_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0875_ (.I(_0034_),
    .Z(net605));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0876_ (.I0(net422),
    .I1(net163),
    .S(_0033_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0877_ (.I(_0035_),
    .Z(net606));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0878_ (.I0(net423),
    .I1(net164),
    .S(_0033_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0879_ (.I(_0036_),
    .Z(net607));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0880_ (.I0(net482),
    .I1(net165),
    .S(_0033_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0881_ (.I(_0037_),
    .Z(net608));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0882_ (.I(_0027_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0883_ (.I0(net489),
    .I1(net166),
    .S(_0038_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0884_ (.I(_0039_),
    .Z(net609));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0885_ (.I0(net490),
    .I1(net167),
    .S(_0038_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0886_ (.I(_0040_),
    .Z(net610));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0887_ (.I0(net492),
    .I1(net168),
    .S(_0038_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0888_ (.I(_0041_),
    .Z(net611));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0889_ (.I0(net493),
    .I1(net169),
    .S(_0038_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0890_ (.I(_0042_),
    .Z(net612));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0891_ (.I(_0027_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0892_ (.I0(net494),
    .I1(net171),
    .S(_0043_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0893_ (.I(_0044_),
    .Z(net614));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0894_ (.I0(net495),
    .I1(net172),
    .S(_0043_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0895_ (.I(_0045_),
    .Z(net615));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0896_ (.I0(net496),
    .I1(net173),
    .S(_0043_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0897_ (.I(_0046_),
    .Z(net616));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0898_ (.I0(net497),
    .I1(net174),
    .S(_0043_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0899_ (.I(_0047_),
    .Z(net617));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0900_ (.I(_0424_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0901_ (.I(_0048_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0902_ (.I0(net498),
    .I1(net175),
    .S(_0049_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0903_ (.I(_0050_),
    .Z(net618));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0904_ (.I0(net483),
    .I1(net176),
    .S(_0049_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0905_ (.I(_0051_),
    .Z(net619));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0906_ (.I0(net484),
    .I1(net177),
    .S(_0049_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0907_ (.I(_0052_),
    .Z(net620));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0908_ (.I0(net485),
    .I1(net178),
    .S(_0049_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0909_ (.I(_0053_),
    .Z(net621));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0910_ (.I(_0048_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0911_ (.I0(net486),
    .I1(net179),
    .S(_0054_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0912_ (.I(_0055_),
    .Z(net622));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0913_ (.I0(net487),
    .I1(net180),
    .S(_0054_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0914_ (.I(_0056_),
    .Z(net623));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0915_ (.I0(net488),
    .I1(net55),
    .S(_0054_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0916_ (.I(_0057_),
    .Z(net499));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0917_ (.I0(_0202_),
    .I1(net56),
    .S(_0054_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0918_ (.I(_0058_),
    .Z(net500));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0919_ (.I(_0048_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0920_ (.I0(_0166_),
    .I1(net57),
    .S(_0059_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0921_ (.I(_0060_),
    .Z(net501));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0922_ (.I0(_0168_),
    .I1(net58),
    .S(_0059_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0923_ (.I(_0061_),
    .Z(net502));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0924_ (.I0(_0164_),
    .I1(net59),
    .S(_0059_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0925_ (.I(_0062_),
    .Z(net503));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0926_ (.I0(_0173_),
    .I1(net60),
    .S(_0059_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0927_ (.I(_0063_),
    .Z(net504));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0928_ (.I(_0048_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0929_ (.I0(_0176_),
    .I1(net61),
    .S(_0064_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0930_ (.I(_0065_),
    .Z(net505));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0931_ (.I0(_0182_),
    .I1(net62),
    .S(_0064_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0932_ (.I(_0066_),
    .Z(net506));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0933_ (.I0(_0186_),
    .I1(net63),
    .S(_0064_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0934_ (.I(_0067_),
    .Z(net507));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0935_ (.I0(_0191_),
    .I1(net64),
    .S(_0064_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0936_ (.I(_0068_),
    .Z(net508));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0937_ (.I(_0424_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0938_ (.I(_0069_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0939_ (.I0(_0194_),
    .I1(net66),
    .S(_0070_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0940_ (.I(_0071_),
    .Z(net510));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0941_ (.I0(_0198_),
    .I1(net67),
    .S(_0070_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0942_ (.I(_0072_),
    .Z(net511));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0943_ (.I0(net699),
    .I1(net68),
    .S(_0070_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0944_ (.I(_0073_),
    .Z(net512));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0945_ (.I0(net698),
    .I1(net69),
    .S(_0070_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0946_ (.I(_0074_),
    .Z(net513));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0947_ (.I(_0069_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0948_ (.I0(net697),
    .I1(net70),
    .S(_0075_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0949_ (.I(_0076_),
    .Z(net514));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0950_ (.I0(net696),
    .I1(net71),
    .S(_0075_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0951_ (.I(_0077_),
    .Z(net515));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0952_ (.I0(net695),
    .I1(net72),
    .S(_0075_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0953_ (.I(_0078_),
    .Z(net516));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0954_ (.I0(net47),
    .I1(net73),
    .S(_0075_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0955_ (.I(_0079_),
    .Z(net517));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0956_ (.I(_0069_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0957_ (.I0(net48),
    .I1(net74),
    .S(_0080_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0958_ (.I(_0081_),
    .Z(net518));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0959_ (.I0(net49),
    .I1(net75),
    .S(_0080_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0960_ (.I(_0082_),
    .Z(net519));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0961_ (.I0(_0265_),
    .I1(net77),
    .S(_0080_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0962_ (.I(_0083_),
    .Z(net521));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0963_ (.A1(_0224_),
    .A2(_0281_),
    .ZN(net473));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0964_ (.I0(net687),
    .I1(net78),
    .S(_0080_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0965_ (.I(_0084_),
    .Z(net522));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0966_ (.I(_0069_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0967_ (.I0(net693),
    .I1(net79),
    .S(_0085_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0968_ (.I(_0086_),
    .Z(net523));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0969_ (.I0(net317),
    .I1(net80),
    .S(_0085_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0970_ (.I(_0087_),
    .Z(net524));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0971_ (.I0(net711),
    .I1(net81),
    .S(_0085_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0972_ (.I(_0088_),
    .Z(net525));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0973_ (.I0(net54),
    .I1(net82),
    .S(_0085_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0974_ (.I(_0089_),
    .Z(net526));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0975_ (.I0(net342),
    .I1(net83),
    .S(_0344_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0976_ (.I(_0090_),
    .Z(net527));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0977_ (.I0(net54),
    .I1(net342),
    .S(_0264_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0978_ (.I(_0091_),
    .Z(net415));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0979_ (.I0(net686),
    .I1(net84),
    .S(_0344_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0980_ (.I(_0092_),
    .Z(net528));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0981_ (.A1(_0203_),
    .A2(_0281_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0982_ (.I(_0093_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0983_ (.I(_0094_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0984_ (.I(_0094_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0985_ (.A1(_0164_),
    .A2(_0096_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0986_ (.A1(_0248_),
    .A2(_0095_),
    .B(_0097_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0987_ (.A1(_0248_),
    .A2(_0250_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0988_ (.I(_0094_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0989_ (.A1(_0173_),
    .A2(_0099_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0990_ (.A1(_0095_),
    .A2(_0098_),
    .B(_0100_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0991_ (.A1(_0248_),
    .A2(_0250_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0992_ (.A1(_0178_),
    .A2(_0101_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0993_ (.A1(_0176_),
    .A2(_0099_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0994_ (.A1(_0095_),
    .A2(_0102_),
    .B(_0103_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0995_ (.A1(\instr_load_addr[0] ),
    .A2(_0250_),
    .A3(_0178_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0996_ (.A1(\instr_load_addr[3] ),
    .A2(_0104_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0997_ (.A1(_0182_),
    .A2(_0099_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0998_ (.A1(_0095_),
    .A2(_0105_),
    .B(_0106_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0999_ (.A1(\instr_load_addr[0] ),
    .A2(\instr_load_addr[1] ),
    .A3(\instr_load_addr[2] ),
    .A4(\instr_load_addr[3] ),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1000_ (.A1(_0187_),
    .A2(_0107_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1001_ (.I(_0093_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1002_ (.I0(_0108_),
    .I1(_0186_),
    .S(_0109_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1003_ (.I(_0110_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1004_ (.A1(_0187_),
    .A2(_0107_),
    .B(\instr_load_addr[5] ),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1005_ (.A1(\instr_load_addr[4] ),
    .A2(\instr_load_addr[5] ),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1006_ (.A1(_0107_),
    .A2(_0112_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1007_ (.I(_0093_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1008_ (.A1(_0191_),
    .A2(_0114_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1009_ (.A1(_0096_),
    .A2(_0111_),
    .A3(_0113_),
    .B(_0115_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1010_ (.I(_0094_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1011_ (.A1(_0195_),
    .A2(_0113_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1012_ (.A1(_0194_),
    .A2(_0099_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1013_ (.A1(_0116_),
    .A2(_0117_),
    .B(_0118_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1014_ (.A1(_0195_),
    .A2(_0113_),
    .B(\instr_load_addr[7] ),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1015_ (.A1(\instr_load_addr[6] ),
    .A2(\instr_load_addr[7] ),
    .A3(_0107_),
    .A4(_0112_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1016_ (.I(_0120_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1017_ (.A1(_0198_),
    .A2(_0109_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1018_ (.A1(_0096_),
    .A2(_0119_),
    .A3(_0121_),
    .B(_0122_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1019_ (.A1(\instr_load_addr[8] ),
    .A2(_0121_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1020_ (.I0(_0123_),
    .I1(net699),
    .S(_0109_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1021_ (.I(_0124_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1022_ (.A1(\instr_load_addr[8] ),
    .A2(_0121_),
    .B(\instr_load_addr[9] ),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1023_ (.A1(\instr_load_addr[8] ),
    .A2(\instr_load_addr[9] ),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1024_ (.A1(_0120_),
    .A2(_0126_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1025_ (.A1(net698),
    .A2(_0109_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1026_ (.A1(_0096_),
    .A2(_0125_),
    .A3(_0127_),
    .B(_0128_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1027_ (.A1(\instr_load_addr[10] ),
    .A2(_0127_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1028_ (.A1(net697),
    .A2(_0114_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1029_ (.A1(_0116_),
    .A2(_0129_),
    .B(_0130_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1030_ (.A1(\instr_load_addr[10] ),
    .A2(_0121_),
    .A3(_0126_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1031_ (.A1(\instr_load_addr[11] ),
    .A2(_0131_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1032_ (.A1(net696),
    .A2(_0114_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1033_ (.A1(_0116_),
    .A2(_0132_),
    .B(_0133_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1034_ (.A1(\instr_load_addr[10] ),
    .A2(\instr_load_addr[11] ),
    .A3(_0120_),
    .A4(_0126_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1035_ (.A1(\instr_load_addr[12] ),
    .A2(_0134_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1036_ (.A1(net695),
    .A2(_0114_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1037_ (.A1(_0116_),
    .A2(_0135_),
    .B(_0136_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1038_ (.A1(_0207_),
    .A2(_0168_),
    .A3(_0281_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1039_ (.I(_0137_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1040_ (.I(_0137_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1041_ (.A1(_0164_),
    .A2(_0139_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1042_ (.A1(_0231_),
    .A2(_0138_),
    .B(_0140_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1043_ (.A1(_0231_),
    .A2(_0235_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1044_ (.A1(_0173_),
    .A2(_0139_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1045_ (.A1(_0138_),
    .A2(_0141_),
    .B(_0142_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1046_ (.A1(_0231_),
    .A2(_0235_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1047_ (.A1(_0177_),
    .A2(_0143_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1048_ (.A1(_0176_),
    .A2(_0139_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1049_ (.A1(_0138_),
    .A2(_0144_),
    .B(_0145_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1050_ (.A1(\data_load_addr[0] ),
    .A2(_0235_),
    .A3(_0177_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1051_ (.A1(\data_load_addr[3] ),
    .A2(_0146_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1052_ (.A1(_0182_),
    .A2(_0139_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1053_ (.A1(_0138_),
    .A2(_0147_),
    .B(_0148_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1054_ (.I(_0137_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1055_ (.A1(\data_load_addr[0] ),
    .A2(\data_load_addr[1] ),
    .A3(\data_load_addr[2] ),
    .A4(\data_load_addr[3] ),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1056_ (.A1(\data_load_addr[4] ),
    .A2(_0150_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1057_ (.A1(\data_load_addr[4] ),
    .A2(_0150_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1058_ (.I(_0137_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1059_ (.A1(_0186_),
    .A2(_0153_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1060_ (.A1(_0149_),
    .A2(_0151_),
    .A3(_0152_),
    .B(_0154_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1061_ (.A1(_0242_),
    .A2(_0151_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1062_ (.A1(_0191_),
    .A2(_0153_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1063_ (.A1(_0149_),
    .A2(_0155_),
    .B(_0156_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1064_ (.A1(_0242_),
    .A2(_0151_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1065_ (.A1(\data_load_addr[6] ),
    .A2(_0157_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1066_ (.A1(_0194_),
    .A2(_0153_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1067_ (.A1(_0149_),
    .A2(_0158_),
    .B(_0159_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1068_ (.A1(_0242_),
    .A2(\data_load_addr[6] ),
    .A3(_0151_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1069_ (.A1(\data_load_addr[7] ),
    .A2(_0160_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1070_ (.A1(_0198_),
    .A2(_0153_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1071_ (.A1(_0149_),
    .A2(_0161_),
    .B(_0162_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1072_ (.A1(net93),
    .A2(net220),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1073_ (.I(_0163_),
    .Z(net643));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1074_ (.D(_0008_),
    .RN(net702),
    .CLK(net678),
    .Q(\instr_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1075_ (.D(_0012_),
    .RN(net700),
    .CLK(net676),
    .Q(\instr_load_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1076_ (.D(_0013_),
    .RN(net700),
    .CLK(net676),
    .Q(\instr_load_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1077_ (.D(_0014_),
    .RN(net700),
    .CLK(net677),
    .Q(\instr_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1078_ (.D(_0015_),
    .RN(net705),
    .CLK(net678),
    .Q(\instr_load_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1079_ (.D(_0016_),
    .RN(net702),
    .CLK(net678),
    .Q(\instr_load_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1080_ (.D(_0017_),
    .RN(net705),
    .CLK(net681),
    .Q(\instr_load_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1081_ (.D(_0018_),
    .RN(net707),
    .CLK(net681),
    .Q(\instr_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1082_ (.D(_0019_),
    .RN(net707),
    .CLK(net681),
    .Q(\instr_load_addr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1083_ (.D(_0020_),
    .RN(net707),
    .CLK(net682),
    .Q(\instr_load_addr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1084_ (.D(_0009_),
    .RN(net708),
    .CLK(net685),
    .Q(\instr_load_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1085_ (.D(_0010_),
    .RN(net708),
    .CLK(net685),
    .Q(\instr_load_addr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1086_ (.D(_0011_),
    .RN(net708),
    .CLK(net685),
    .Q(\instr_load_addr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1087_ (.D(_0000_),
    .RN(net700),
    .CLK(net676),
    .Q(\data_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1088_ (.D(_0001_),
    .RN(net701),
    .CLK(net676),
    .Q(\data_load_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1089_ (.D(_0002_),
    .RN(net701),
    .CLK(net677),
    .Q(\data_load_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1090_ (.D(_0003_),
    .RN(net703),
    .CLK(net677),
    .Q(\data_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1091_ (.D(_0004_),
    .RN(net703),
    .CLK(net678),
    .Q(\data_load_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1092_ (.D(_0005_),
    .RN(net705),
    .CLK(net679),
    .Q(\data_load_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1093_ (.D(_0006_),
    .RN(net706),
    .CLK(net681),
    .Q(\data_load_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1094_ (.D(_0007_),
    .RN(net707),
    .CLK(net682),
    .Q(\data_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_759 (.Z(net759));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_760 (.Z(net760));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_761 (.Z(net761));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_762 (.Z(net762));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_763 (.Z(net763));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_764 (.Z(net764));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_765 (.Z(net765));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_766 (.Z(net766));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_767 (.Z(net767));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_768 (.Z(net768));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_769 (.Z(net769));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_770 (.Z(net770));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_771 (.Z(net771));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_772 (.Z(net772));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_773 (.Z(net773));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_774 (.Z(net774));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_775 (.Z(net775));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_776 (.Z(net776));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_777 (.Z(net777));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_778 (.Z(net778));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0891__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_713 (.ZN(net713));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_714 (.ZN(net714));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_715 (.ZN(net715));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_716 (.ZN(net716));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_717 (.ZN(net717));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_718 (.ZN(net718));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_719 (.ZN(net719));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_720 (.ZN(net720));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_721 (.ZN(net721));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_722 (.ZN(net722));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_723 (.ZN(net723));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_724 (.ZN(net724));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_725 (.ZN(net725));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_726 (.ZN(net726));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_727 (.ZN(net727));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_728 (.ZN(net728));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_729 (.ZN(net729));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_730 (.ZN(net730));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_731 (.ZN(net731));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_732 (.ZN(net732));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_733 (.ZN(net733));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_734 (.ZN(net734));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_735 (.ZN(net735));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_736 (.ZN(net736));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_737 (.ZN(net737));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_738 (.ZN(net738));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_739 (.ZN(net739));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_740 (.ZN(net740));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_741 (.ZN(net741));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_742 (.ZN(net742));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_743 (.ZN(net743));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_744 (.ZN(net744));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_745 (.ZN(net745));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_746 (.ZN(net746));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_747 (.ZN(net747));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_748 (.ZN(net748));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_749 (.ZN(net749));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_750 (.ZN(net750));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_751 (.ZN(net751));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_752 (.ZN(net752));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_753 (.ZN(net753));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_754 (.ZN(net754));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_755 (.ZN(net755));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_756 (.ZN(net756));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_757 (.ZN(net757));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_758 (.Z(net758));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1162_ (.I(net344),
    .Z(analog_io[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1163_ (.I(net355),
    .Z(analog_io[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1164_ (.I(net366),
    .Z(analog_io[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1165_ (.I(net369),
    .Z(analog_io[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1166_ (.I(net370),
    .Z(analog_io[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1167_ (.I(net371),
    .Z(analog_io[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1168_ (.I(net372),
    .Z(analog_io[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1169_ (.I(net373),
    .Z(analog_io[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1170_ (.I(net374),
    .Z(analog_io[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1171_ (.I(net375),
    .Z(analog_io[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1172_ (.I(net345),
    .Z(analog_io[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1173_ (.I(net346),
    .Z(analog_io[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1174_ (.I(net347),
    .Z(analog_io[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1175_ (.I(net348),
    .Z(analog_io[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1176_ (.I(net349),
    .Z(analog_io[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1177_ (.I(net350),
    .Z(analog_io[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1178_ (.I(net351),
    .Z(analog_io[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1179_ (.I(net352),
    .Z(analog_io[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1180_ (.I(net353),
    .Z(analog_io[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1181_ (.I(net354),
    .Z(analog_io[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1182_ (.I(net356),
    .Z(analog_io[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1183_ (.I(net357),
    .Z(analog_io[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1184_ (.I(net358),
    .Z(analog_io[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1185_ (.I(net359),
    .Z(analog_io[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1186_ (.I(net360),
    .Z(analog_io[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1187_ (.I(net361),
    .Z(analog_io[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1188_ (.I(net362),
    .Z(analog_io[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1189_ (.I(net363),
    .Z(analog_io[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1190_ (.I(net364),
    .Z(analog_io[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1191_ (.I(net691),
    .Z(net441));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1192_ (.I(net691),
    .Z(net442));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1193_ (.I(net691),
    .Z(net443));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1194_ (.I(net692),
    .Z(net444));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1195_ (.I(net692),
    .Z(net445));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1196_ (.I(net692),
    .Z(net446));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1197_ (.I(net693),
    .Z(net447));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1198_ (.I(net440),
    .Z(net448));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1199_ (.I(net34),
    .Z(net457));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1200_ (.I(net35),
    .Z(net464));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1201_ (.I(net36),
    .Z(net465));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1202_ (.I(net37),
    .Z(net466));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1203_ (.I(net38),
    .Z(net467));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1204_ (.I(net39),
    .Z(net468));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1205_ (.I(net40),
    .Z(net469));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1206_ (.I(net41),
    .Z(net470));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1207_ (.I(net42),
    .Z(net471));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1208_ (.I(net43),
    .Z(net472));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1209_ (.I(net44),
    .Z(net458));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1210_ (.I(net45),
    .Z(net459));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1211_ (.I(net46),
    .Z(net460));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1212_ (.I(net47),
    .Z(net461));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1213_ (.I(net48),
    .Z(net462));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1214_ (.I(net49),
    .Z(net463));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1215_ (.I(net690),
    .Z(net474));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1216_ (.I(net690),
    .Z(net475));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1217_ (.I(net689),
    .Z(net476));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1218_ (.I(net688),
    .Z(net477));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1219_ (.I(net687),
    .Z(net478));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1220_ (.I(net687),
    .Z(net479));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1221_ (.I(net687),
    .Z(net480));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1222_ (.I(net688),
    .Z(net481));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1223_ (.I(net17),
    .Z(net491));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1224_ (.I(net711),
    .Z(net625));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1225_ (.I(net53),
    .Z(net626));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1226_ (.I(net377),
    .Z(net644));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1227_ (.I(net388),
    .Z(net655));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1228_ (.I(net399),
    .Z(net666));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1229_ (.I(net402),
    .Z(net669));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1230_ (.I(net403),
    .Z(net670));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1231_ (.I(net404),
    .Z(net671));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1232_ (.I(net405),
    .Z(net672));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1233_ (.I(net406),
    .Z(net673));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1234_ (.I(net407),
    .Z(net674));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1235_ (.I(net408),
    .Z(net675));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1236_ (.I(net378),
    .Z(net645));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1237_ (.I(net379),
    .Z(net646));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1238_ (.I(net380),
    .Z(net647));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1239_ (.I(net381),
    .Z(net648));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1240_ (.I(net382),
    .Z(net649));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1241_ (.I(net383),
    .Z(net650));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1242_ (.I(net384),
    .Z(net651));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1243_ (.I(net385),
    .Z(net652));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1244_ (.I(net386),
    .Z(net653));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1245_ (.I(net387),
    .Z(net654));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1246_ (.I(net389),
    .Z(net656));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1247_ (.I(net390),
    .Z(net657));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1248_ (.I(net391),
    .Z(net658));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1249_ (.I(net392),
    .Z(net659));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1250_ (.I(net393),
    .Z(net660));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1251_ (.I(net394),
    .Z(net661));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1252_ (.I(net395),
    .Z(net662));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1253_ (.I(net396),
    .Z(net663));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1254_ (.I(net397),
    .Z(net664));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1255_ (.I(net398),
    .Z(net665));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1256_ (.I(net400),
    .Z(net667));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1257_ (.I(net401),
    .Z(net668));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11577 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(data_read_data[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(data_read_data[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(data_read_data[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(data_read_data[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(data_read_data[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(data_read_data[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input7 (.I(data_read_data[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(data_read_data[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(data_read_data[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(data_read_data[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(data_read_data[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(data_read_data[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(data_read_data[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(data_read_data[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input15 (.I(data_read_data[8]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(data_read_data[9]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input17 (.I(hlt),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(instr[0]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(instr[10]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(instr[11]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(instr[12]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input22 (.I(instr[13]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input23 (.I(instr[14]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input24 (.I(instr[15]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(instr[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(instr[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input27 (.I(instr[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(instr[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input29 (.I(instr[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input30 (.I(instr[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(instr[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(instr[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(instr[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input34 (.I(io_in[16]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input35 (.I(io_in[17]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(io_in[18]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input37 (.I(io_in[19]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input38 (.I(io_in[20]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input39 (.I(io_in[21]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(io_in[22]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input41 (.I(io_in[23]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(io_in[24]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(io_in[25]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(io_in[26]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(io_in[27]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input46 (.I(io_in[28]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input47 (.I(io_in[29]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input48 (.I(io_in[30]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input49 (.I(io_in[31]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input50 (.I(io_in[32]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(io_in[33]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input52 (.I(io_in[34]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input53 (.I(io_in[36]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input54 (.I(io_in[37]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input55 (.I(la_data_in[100]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input56 (.I(la_data_in[101]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input57 (.I(la_data_in[102]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input58 (.I(la_data_in[103]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input59 (.I(la_data_in[104]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input60 (.I(la_data_in[105]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input61 (.I(la_data_in[106]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input62 (.I(la_data_in[107]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input63 (.I(la_data_in[108]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input64 (.I(la_data_in[109]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input65 (.I(la_data_in[10]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input66 (.I(la_data_in[110]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input67 (.I(la_data_in[111]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input68 (.I(la_data_in[112]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input69 (.I(la_data_in[113]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input70 (.I(la_data_in[114]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input71 (.I(la_data_in[115]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input72 (.I(la_data_in[116]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input73 (.I(la_data_in[117]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input74 (.I(la_data_in[118]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input75 (.I(la_data_in[119]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input76 (.I(la_data_in[11]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input77 (.I(la_data_in[120]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input78 (.I(la_data_in[121]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input79 (.I(la_data_in[122]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input80 (.I(la_data_in[123]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input81 (.I(la_data_in[124]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input82 (.I(la_data_in[125]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input83 (.I(la_data_in[126]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input84 (.I(la_data_in[127]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input85 (.I(la_data_in[12]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input86 (.I(la_data_in[13]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input87 (.I(la_data_in[14]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input88 (.I(la_data_in[15]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input89 (.I(la_data_in[16]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input90 (.I(la_data_in[17]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input91 (.I(la_data_in[18]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input92 (.I(la_data_in[19]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input93 (.I(la_data_in[1]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input94 (.I(la_data_in[20]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input95 (.I(la_data_in[21]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input96 (.I(la_data_in[22]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input97 (.I(la_data_in[23]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input98 (.I(la_data_in[24]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input99 (.I(la_data_in[25]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input100 (.I(la_data_in[26]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input101 (.I(la_data_in[27]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input102 (.I(la_data_in[28]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input103 (.I(la_data_in[29]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input104 (.I(la_data_in[2]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input105 (.I(la_data_in[30]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input106 (.I(la_data_in[31]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input107 (.I(la_data_in[32]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input108 (.I(la_data_in[33]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input109 (.I(la_data_in[34]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input110 (.I(la_data_in[35]),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input111 (.I(la_data_in[36]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input112 (.I(la_data_in[37]),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input113 (.I(la_data_in[38]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input114 (.I(la_data_in[39]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input115 (.I(la_data_in[3]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input116 (.I(la_data_in[40]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input117 (.I(la_data_in[41]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input118 (.I(la_data_in[42]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input119 (.I(la_data_in[43]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input120 (.I(la_data_in[44]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input121 (.I(la_data_in[45]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input122 (.I(la_data_in[46]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input123 (.I(la_data_in[47]),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input124 (.I(la_data_in[48]),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input125 (.I(la_data_in[49]),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input126 (.I(la_data_in[4]),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input127 (.I(la_data_in[50]),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input128 (.I(la_data_in[51]),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input129 (.I(la_data_in[52]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input130 (.I(la_data_in[53]),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input131 (.I(la_data_in[54]),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input132 (.I(la_data_in[55]),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input133 (.I(la_data_in[56]),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input134 (.I(la_data_in[57]),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input135 (.I(la_data_in[58]),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input136 (.I(la_data_in[59]),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input137 (.I(la_data_in[5]),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input138 (.I(la_data_in[60]),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input139 (.I(la_data_in[61]),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input140 (.I(la_data_in[62]),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input141 (.I(la_data_in[63]),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input142 (.I(la_data_in[64]),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input143 (.I(la_data_in[65]),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input144 (.I(la_data_in[66]),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input145 (.I(la_data_in[67]),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input146 (.I(la_data_in[68]),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input147 (.I(la_data_in[69]),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input148 (.I(la_data_in[6]),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input149 (.I(la_data_in[70]),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input150 (.I(la_data_in[71]),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input151 (.I(la_data_in[72]),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input152 (.I(la_data_in[73]),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input153 (.I(la_data_in[74]),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input154 (.I(la_data_in[75]),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input155 (.I(la_data_in[76]),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input156 (.I(la_data_in[77]),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input157 (.I(la_data_in[78]),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input158 (.I(la_data_in[79]),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input159 (.I(la_data_in[7]),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input160 (.I(la_data_in[80]),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input161 (.I(la_data_in[81]),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input162 (.I(la_data_in[82]),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input163 (.I(la_data_in[83]),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input164 (.I(la_data_in[84]),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input165 (.I(la_data_in[85]),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input166 (.I(la_data_in[86]),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input167 (.I(la_data_in[87]),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input168 (.I(la_data_in[88]),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input169 (.I(la_data_in[89]),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input170 (.I(la_data_in[8]),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input171 (.I(la_data_in[90]),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input172 (.I(la_data_in[91]),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input173 (.I(la_data_in[92]),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input174 (.I(la_data_in[93]),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input175 (.I(la_data_in[94]),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input176 (.I(la_data_in[95]),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input177 (.I(la_data_in[96]),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input178 (.I(la_data_in[97]),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input179 (.I(la_data_in[98]),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input180 (.I(la_data_in[99]),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input181 (.I(la_data_in[9]),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input182 (.I(la_oenb[100]),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input183 (.I(la_oenb[101]),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input184 (.I(la_oenb[102]),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input185 (.I(la_oenb[103]),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input186 (.I(la_oenb[104]),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input187 (.I(la_oenb[105]),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input188 (.I(la_oenb[106]),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input189 (.I(la_oenb[107]),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input190 (.I(la_oenb[108]),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input191 (.I(la_oenb[109]),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input192 (.I(la_oenb[10]),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input193 (.I(la_oenb[110]),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input194 (.I(la_oenb[111]),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input195 (.I(la_oenb[112]),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input196 (.I(la_oenb[113]),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input197 (.I(la_oenb[114]),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input198 (.I(la_oenb[115]),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input199 (.I(la_oenb[116]),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input200 (.I(la_oenb[117]),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input201 (.I(la_oenb[118]),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input202 (.I(la_oenb[119]),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input203 (.I(la_oenb[11]),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input204 (.I(la_oenb[120]),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input205 (.I(la_oenb[121]),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input206 (.I(la_oenb[122]),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input207 (.I(la_oenb[123]),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input208 (.I(la_oenb[124]),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input209 (.I(la_oenb[125]),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input210 (.I(la_oenb[126]),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input211 (.I(la_oenb[127]),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input212 (.I(la_oenb[12]),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input213 (.I(la_oenb[13]),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input214 (.I(la_oenb[14]),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input215 (.I(la_oenb[15]),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input216 (.I(la_oenb[16]),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input217 (.I(la_oenb[17]),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input218 (.I(la_oenb[18]),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input219 (.I(la_oenb[19]),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input220 (.I(la_oenb[1]),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input221 (.I(la_oenb[20]),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input222 (.I(la_oenb[21]),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input223 (.I(la_oenb[22]),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input224 (.I(la_oenb[23]),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input225 (.I(la_oenb[24]),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input226 (.I(la_oenb[25]),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input227 (.I(la_oenb[26]),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input228 (.I(la_oenb[27]),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input229 (.I(la_oenb[28]),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input230 (.I(la_oenb[29]),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input231 (.I(la_oenb[2]),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input232 (.I(la_oenb[30]),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input233 (.I(la_oenb[31]),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input234 (.I(la_oenb[32]),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input235 (.I(la_oenb[33]),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input236 (.I(la_oenb[34]),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input237 (.I(la_oenb[35]),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input238 (.I(la_oenb[36]),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input239 (.I(la_oenb[37]),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input240 (.I(la_oenb[38]),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input241 (.I(la_oenb[39]),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input242 (.I(la_oenb[3]),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input243 (.I(la_oenb[40]),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input244 (.I(la_oenb[41]),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input245 (.I(la_oenb[42]),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input246 (.I(la_oenb[43]),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input247 (.I(la_oenb[44]),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input248 (.I(la_oenb[45]),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input249 (.I(la_oenb[46]),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input250 (.I(la_oenb[47]),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input251 (.I(la_oenb[48]),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input252 (.I(la_oenb[49]),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input253 (.I(la_oenb[4]),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input254 (.I(la_oenb[50]),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input255 (.I(la_oenb[51]),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input256 (.I(la_oenb[52]),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input257 (.I(la_oenb[53]),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input258 (.I(la_oenb[54]),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input259 (.I(la_oenb[55]),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input260 (.I(la_oenb[56]),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input261 (.I(la_oenb[57]),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input262 (.I(la_oenb[58]),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input263 (.I(la_oenb[59]),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input264 (.I(la_oenb[5]),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input265 (.I(la_oenb[60]),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input266 (.I(la_oenb[61]),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input267 (.I(la_oenb[62]),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input268 (.I(la_oenb[63]),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input269 (.I(la_oenb[64]),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input270 (.I(la_oenb[65]),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input271 (.I(la_oenb[66]),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input272 (.I(la_oenb[67]),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input273 (.I(la_oenb[68]),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input274 (.I(la_oenb[69]),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input275 (.I(la_oenb[6]),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input276 (.I(la_oenb[70]),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input277 (.I(la_oenb[71]),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input278 (.I(la_oenb[72]),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input279 (.I(la_oenb[73]),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input280 (.I(la_oenb[74]),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input281 (.I(la_oenb[75]),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input282 (.I(la_oenb[76]),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input283 (.I(la_oenb[77]),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input284 (.I(la_oenb[78]),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input285 (.I(la_oenb[79]),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input286 (.I(la_oenb[7]),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input287 (.I(la_oenb[80]),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input288 (.I(la_oenb[81]),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input289 (.I(la_oenb[82]),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input290 (.I(la_oenb[83]),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input291 (.I(la_oenb[84]),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input292 (.I(la_oenb[85]),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input293 (.I(la_oenb[86]),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input294 (.I(la_oenb[87]),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input295 (.I(la_oenb[88]),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input296 (.I(la_oenb[89]),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input297 (.I(la_oenb[8]),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input298 (.I(la_oenb[90]),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input299 (.I(la_oenb[91]),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input300 (.I(la_oenb[92]),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input301 (.I(la_oenb[93]),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input302 (.I(la_oenb[94]),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input303 (.I(la_oenb[95]),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input304 (.I(la_oenb[96]),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input305 (.I(la_oenb[97]),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input306 (.I(la_oenb[98]),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input307 (.I(la_oenb[99]),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input308 (.I(la_oenb[9]),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input309 (.I(uP_data_mem_addr[0]),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input310 (.I(uP_data_mem_addr[1]),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input311 (.I(uP_data_mem_addr[2]),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input312 (.I(uP_data_mem_addr[3]),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input313 (.I(uP_data_mem_addr[4]),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input314 (.I(uP_data_mem_addr[5]),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input315 (.I(uP_data_mem_addr[6]),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input316 (.I(uP_data_mem_addr[7]),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input317 (.I(uP_dataw_en),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input318 (.I(uP_instr_mem_addr[0]),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input319 (.I(uP_instr_mem_addr[1]),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input320 (.I(uP_instr_mem_addr[2]),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input321 (.I(uP_instr_mem_addr[3]),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input322 (.I(uP_instr_mem_addr[4]),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input323 (.I(uP_instr_mem_addr[5]),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input324 (.I(uP_instr_mem_addr[6]),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input325 (.I(uP_instr_mem_addr[7]),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input326 (.I(uP_write_data[0]),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input327 (.I(uP_write_data[10]),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input328 (.I(uP_write_data[11]),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input329 (.I(uP_write_data[12]),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input330 (.I(uP_write_data[13]),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input331 (.I(uP_write_data[14]),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input332 (.I(uP_write_data[15]),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input333 (.I(uP_write_data[1]),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input334 (.I(uP_write_data[2]),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input335 (.I(uP_write_data[3]),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input336 (.I(uP_write_data[4]),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input337 (.I(uP_write_data[5]),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input338 (.I(uP_write_data[6]),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input339 (.I(uP_write_data[7]),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input340 (.I(uP_write_data[8]),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input341 (.I(uP_write_data[9]),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input342 (.I(wb_clk_i),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input343 (.I(wb_rst_i),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input344 (.I(wbs_adr_i[0]),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input345 (.I(wbs_adr_i[10]),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input346 (.I(wbs_adr_i[11]),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input347 (.I(wbs_adr_i[12]),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input348 (.I(wbs_adr_i[13]),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input349 (.I(wbs_adr_i[14]),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input350 (.I(wbs_adr_i[15]),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input351 (.I(wbs_adr_i[16]),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input352 (.I(wbs_adr_i[17]),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input353 (.I(wbs_adr_i[18]),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input354 (.I(wbs_adr_i[19]),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input355 (.I(wbs_adr_i[1]),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input356 (.I(wbs_adr_i[20]),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input357 (.I(wbs_adr_i[21]),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input358 (.I(wbs_adr_i[22]),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input359 (.I(wbs_adr_i[23]),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input360 (.I(wbs_adr_i[24]),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input361 (.I(wbs_adr_i[25]),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input362 (.I(wbs_adr_i[26]),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input363 (.I(wbs_adr_i[27]),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input364 (.I(wbs_adr_i[28]),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input365 (.I(wbs_adr_i[29]),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input366 (.I(wbs_adr_i[2]),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input367 (.I(wbs_adr_i[30]),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input368 (.I(wbs_adr_i[31]),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input369 (.I(wbs_adr_i[3]),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input370 (.I(wbs_adr_i[4]),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input371 (.I(wbs_adr_i[5]),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input372 (.I(wbs_adr_i[6]),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input373 (.I(wbs_adr_i[7]),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input374 (.I(wbs_adr_i[8]),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input375 (.I(wbs_adr_i[9]),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input376 (.I(wbs_cyc_i),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input377 (.I(wbs_dat_i[0]),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input378 (.I(wbs_dat_i[10]),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input379 (.I(wbs_dat_i[11]),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input380 (.I(wbs_dat_i[12]),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input381 (.I(wbs_dat_i[13]),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input382 (.I(wbs_dat_i[14]),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input383 (.I(wbs_dat_i[15]),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input384 (.I(wbs_dat_i[16]),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input385 (.I(wbs_dat_i[17]),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input386 (.I(wbs_dat_i[18]),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input387 (.I(wbs_dat_i[19]),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input388 (.I(wbs_dat_i[1]),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input389 (.I(wbs_dat_i[20]),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input390 (.I(wbs_dat_i[21]),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input391 (.I(wbs_dat_i[22]),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input392 (.I(wbs_dat_i[23]),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input393 (.I(wbs_dat_i[24]),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input394 (.I(wbs_dat_i[25]),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input395 (.I(wbs_dat_i[26]),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input396 (.I(wbs_dat_i[27]),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input397 (.I(wbs_dat_i[28]),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input398 (.I(wbs_dat_i[29]),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input399 (.I(wbs_dat_i[2]),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input400 (.I(wbs_dat_i[30]),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input401 (.I(wbs_dat_i[31]),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input402 (.I(wbs_dat_i[3]),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input403 (.I(wbs_dat_i[4]),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input404 (.I(wbs_dat_i[5]),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input405 (.I(wbs_dat_i[6]),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input406 (.I(wbs_dat_i[7]),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input407 (.I(wbs_dat_i[8]),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input408 (.I(wbs_dat_i[9]),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input409 (.I(wbs_sel_i[0]),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input410 (.I(wbs_sel_i[1]),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input411 (.I(wbs_sel_i[2]),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input412 (.I(wbs_sel_i[3]),
    .Z(net412));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input413 (.I(wbs_stb_i),
    .Z(net413));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input414 (.I(wbs_we_i),
    .Z(net414));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output415 (.I(net686),
    .Z(clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output416 (.I(net416),
    .Z(data_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output417 (.I(net417),
    .Z(data_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output418 (.I(net418),
    .Z(data_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output419 (.I(net419),
    .Z(data_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output420 (.I(net420),
    .Z(data_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output421 (.I(net421),
    .Z(data_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output422 (.I(net422),
    .Z(data_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output423 (.I(net423),
    .Z(data_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output424 (.I(net424),
    .Z(data_write_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output425 (.I(net425),
    .Z(data_write_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output426 (.I(net426),
    .Z(data_write_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output427 (.I(net427),
    .Z(data_write_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output428 (.I(net428),
    .Z(data_write_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output429 (.I(net429),
    .Z(data_write_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output430 (.I(net430),
    .Z(data_write_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output431 (.I(net431),
    .Z(data_write_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output432 (.I(net432),
    .Z(data_write_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output433 (.I(net433),
    .Z(data_write_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output434 (.I(net434),
    .Z(data_write_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output435 (.I(net435),
    .Z(data_write_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output436 (.I(net436),
    .Z(data_write_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output437 (.I(net437),
    .Z(data_write_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output438 (.I(net438),
    .Z(data_write_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output439 (.I(net439),
    .Z(data_write_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output440 (.I(net691),
    .Z(dataw_en));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output441 (.I(net441),
    .Z(dataw_en_8bit[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output442 (.I(net442),
    .Z(dataw_en_8bit[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output443 (.I(net443),
    .Z(dataw_en_8bit[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output444 (.I(net444),
    .Z(dataw_en_8bit[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output445 (.I(net445),
    .Z(dataw_en_8bit[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output446 (.I(net446),
    .Z(dataw_en_8bit[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output447 (.I(net447),
    .Z(dataw_en_8bit[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output448 (.I(net448),
    .Z(dataw_en_8bit[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output449 (.I(net449),
    .Z(instr_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output450 (.I(net450),
    .Z(instr_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output451 (.I(net451),
    .Z(instr_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output452 (.I(net452),
    .Z(instr_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output453 (.I(net453),
    .Z(instr_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output454 (.I(net454),
    .Z(instr_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output455 (.I(net455),
    .Z(instr_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output456 (.I(net456),
    .Z(instr_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output457 (.I(net457),
    .Z(instr_write_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output458 (.I(net458),
    .Z(instr_write_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output459 (.I(net459),
    .Z(instr_write_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output460 (.I(net460),
    .Z(instr_write_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output461 (.I(net461),
    .Z(instr_write_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output462 (.I(net462),
    .Z(instr_write_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output463 (.I(net463),
    .Z(instr_write_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output464 (.I(net464),
    .Z(instr_write_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output465 (.I(net465),
    .Z(instr_write_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output466 (.I(net466),
    .Z(instr_write_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output467 (.I(net467),
    .Z(instr_write_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output468 (.I(net468),
    .Z(instr_write_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output469 (.I(net469),
    .Z(instr_write_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output470 (.I(net470),
    .Z(instr_write_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output471 (.I(net471),
    .Z(instr_write_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output472 (.I(net472),
    .Z(instr_write_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output473 (.I(net690),
    .Z(instrw_en));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output474 (.I(net474),
    .Z(instrw_en_8bit[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output475 (.I(net475),
    .Z(instrw_en_8bit[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output476 (.I(net476),
    .Z(instrw_en_8bit[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output477 (.I(net477),
    .Z(instrw_en_8bit[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output478 (.I(net478),
    .Z(instrw_en_8bit[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output479 (.I(net479),
    .Z(instrw_en_8bit[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output480 (.I(net480),
    .Z(instrw_en_8bit[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output481 (.I(net481),
    .Z(instrw_en_8bit[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output482 (.I(net482),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output483 (.I(net483),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output484 (.I(net484),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output485 (.I(net485),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output486 (.I(net486),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output487 (.I(net487),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output488 (.I(net488),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output489 (.I(net489),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output490 (.I(net490),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output491 (.I(net491),
    .Z(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output492 (.I(net492),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output493 (.I(net493),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output494 (.I(net494),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output495 (.I(net495),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output496 (.I(net496),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output497 (.I(net497),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output498 (.I(net498),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output499 (.I(net499),
    .Z(la_data_out[100]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output500 (.I(net500),
    .Z(la_data_out[101]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output501 (.I(net501),
    .Z(la_data_out[102]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output502 (.I(net502),
    .Z(la_data_out[103]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output503 (.I(net503),
    .Z(la_data_out[104]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output504 (.I(net504),
    .Z(la_data_out[105]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output505 (.I(net505),
    .Z(la_data_out[106]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output506 (.I(net506),
    .Z(la_data_out[107]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output507 (.I(net507),
    .Z(la_data_out[108]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output508 (.I(net508),
    .Z(la_data_out[109]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output509 (.I(net509),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output510 (.I(net510),
    .Z(la_data_out[110]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output511 (.I(net511),
    .Z(la_data_out[111]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output512 (.I(net512),
    .Z(la_data_out[112]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output513 (.I(net513),
    .Z(la_data_out[113]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output514 (.I(net514),
    .Z(la_data_out[114]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output515 (.I(net515),
    .Z(la_data_out[115]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output516 (.I(net516),
    .Z(la_data_out[116]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output517 (.I(net517),
    .Z(la_data_out[117]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output518 (.I(net518),
    .Z(la_data_out[118]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output519 (.I(net519),
    .Z(la_data_out[119]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output520 (.I(net520),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output521 (.I(net521),
    .Z(la_data_out[120]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output522 (.I(net522),
    .Z(la_data_out[121]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output523 (.I(net523),
    .Z(la_data_out[122]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output524 (.I(net524),
    .Z(la_data_out[123]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output525 (.I(net525),
    .Z(la_data_out[124]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output526 (.I(net526),
    .Z(la_data_out[125]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output527 (.I(net527),
    .Z(la_data_out[126]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output528 (.I(net528),
    .Z(la_data_out[127]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output529 (.I(net529),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output530 (.I(net530),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output531 (.I(net531),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output532 (.I(net532),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output533 (.I(net533),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output534 (.I(net534),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output535 (.I(net535),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output536 (.I(net536),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output537 (.I(net537),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output538 (.I(net538),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output539 (.I(net539),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output540 (.I(net540),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output541 (.I(net541),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output542 (.I(net542),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output543 (.I(net543),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output544 (.I(net544),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output545 (.I(net545),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output546 (.I(net546),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output547 (.I(net547),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output548 (.I(net548),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output549 (.I(net549),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output550 (.I(net550),
    .Z(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output551 (.I(net551),
    .Z(la_data_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output552 (.I(net552),
    .Z(la_data_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output553 (.I(net553),
    .Z(la_data_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output554 (.I(net554),
    .Z(la_data_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output555 (.I(net555),
    .Z(la_data_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output556 (.I(net556),
    .Z(la_data_out[38]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output557 (.I(net557),
    .Z(la_data_out[39]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output558 (.I(net558),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output559 (.I(net559),
    .Z(la_data_out[40]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output560 (.I(net560),
    .Z(la_data_out[41]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output561 (.I(net561),
    .Z(la_data_out[42]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output562 (.I(net562),
    .Z(la_data_out[43]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output563 (.I(net563),
    .Z(la_data_out[44]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output564 (.I(net564),
    .Z(la_data_out[45]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output565 (.I(net565),
    .Z(la_data_out[46]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output566 (.I(net566),
    .Z(la_data_out[47]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output567 (.I(net567),
    .Z(la_data_out[48]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output568 (.I(net568),
    .Z(la_data_out[49]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output569 (.I(net569),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output570 (.I(net570),
    .Z(la_data_out[50]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output571 (.I(net571),
    .Z(la_data_out[51]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output572 (.I(net572),
    .Z(la_data_out[52]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output573 (.I(net573),
    .Z(la_data_out[53]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output574 (.I(net574),
    .Z(la_data_out[54]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output575 (.I(net575),
    .Z(la_data_out[55]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output576 (.I(net576),
    .Z(la_data_out[56]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output577 (.I(net577),
    .Z(la_data_out[57]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output578 (.I(net578),
    .Z(la_data_out[58]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output579 (.I(net579),
    .Z(la_data_out[59]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output580 (.I(net580),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output581 (.I(net581),
    .Z(la_data_out[60]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output582 (.I(net582),
    .Z(la_data_out[61]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output583 (.I(net583),
    .Z(la_data_out[62]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output584 (.I(net584),
    .Z(la_data_out[63]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output585 (.I(net585),
    .Z(la_data_out[64]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output586 (.I(net586),
    .Z(la_data_out[65]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output587 (.I(net587),
    .Z(la_data_out[66]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output588 (.I(net588),
    .Z(la_data_out[67]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output589 (.I(net589),
    .Z(la_data_out[68]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output590 (.I(net590),
    .Z(la_data_out[69]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output591 (.I(net591),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output592 (.I(net592),
    .Z(la_data_out[70]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output593 (.I(net593),
    .Z(la_data_out[71]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output594 (.I(net594),
    .Z(la_data_out[72]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output595 (.I(net595),
    .Z(la_data_out[73]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output596 (.I(net596),
    .Z(la_data_out[74]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output597 (.I(net597),
    .Z(la_data_out[75]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output598 (.I(net598),
    .Z(la_data_out[76]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output599 (.I(net599),
    .Z(la_data_out[77]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output600 (.I(net600),
    .Z(la_data_out[78]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output601 (.I(net601),
    .Z(la_data_out[79]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output602 (.I(net602),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output603 (.I(net603),
    .Z(la_data_out[80]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output604 (.I(net604),
    .Z(la_data_out[81]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output605 (.I(net605),
    .Z(la_data_out[82]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output606 (.I(net606),
    .Z(la_data_out[83]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output607 (.I(net607),
    .Z(la_data_out[84]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output608 (.I(net608),
    .Z(la_data_out[85]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output609 (.I(net609),
    .Z(la_data_out[86]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output610 (.I(net610),
    .Z(la_data_out[87]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output611 (.I(net611),
    .Z(la_data_out[88]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output612 (.I(net612),
    .Z(la_data_out[89]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output613 (.I(net613),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output614 (.I(net614),
    .Z(la_data_out[90]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output615 (.I(net615),
    .Z(la_data_out[91]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output616 (.I(net616),
    .Z(la_data_out[92]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output617 (.I(net617),
    .Z(la_data_out[93]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output618 (.I(net618),
    .Z(la_data_out[94]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output619 (.I(net619),
    .Z(la_data_out[95]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output620 (.I(net620),
    .Z(la_data_out[96]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output621 (.I(net621),
    .Z(la_data_out[97]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output622 (.I(net622),
    .Z(la_data_out[98]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output623 (.I(net623),
    .Z(la_data_out[99]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output624 (.I(net624),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output625 (.I(net625),
    .Z(reset));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output626 (.I(net626),
    .Z(start));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output627 (.I(net627),
    .Z(uP_instr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output628 (.I(net628),
    .Z(uP_instr[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output629 (.I(net629),
    .Z(uP_instr[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output630 (.I(net630),
    .Z(uP_instr[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output631 (.I(net631),
    .Z(uP_instr[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output632 (.I(net632),
    .Z(uP_instr[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output633 (.I(net633),
    .Z(uP_instr[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output634 (.I(net634),
    .Z(uP_instr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output635 (.I(net635),
    .Z(uP_instr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output636 (.I(net636),
    .Z(uP_instr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output637 (.I(net637),
    .Z(uP_instr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output638 (.I(net638),
    .Z(uP_instr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output639 (.I(net639),
    .Z(uP_instr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output640 (.I(net640),
    .Z(uP_instr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output641 (.I(net641),
    .Z(uP_instr[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output642 (.I(net642),
    .Z(uP_instr[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output643 (.I(net643),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output644 (.I(net644),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output645 (.I(net645),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output646 (.I(net646),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output647 (.I(net647),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output648 (.I(net648),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output649 (.I(net649),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output650 (.I(net650),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output651 (.I(net651),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output652 (.I(net652),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output653 (.I(net653),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output654 (.I(net654),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output655 (.I(net655),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output656 (.I(net656),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output657 (.I(net657),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output658 (.I(net658),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output659 (.I(net659),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output660 (.I(net660),
    .Z(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output661 (.I(net661),
    .Z(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output662 (.I(net662),
    .Z(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output663 (.I(net663),
    .Z(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output664 (.I(net664),
    .Z(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output665 (.I(net665),
    .Z(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output666 (.I(net666),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output667 (.I(net667),
    .Z(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output668 (.I(net668),
    .Z(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output669 (.I(net669),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output670 (.I(net670),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output671 (.I(net671),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output672 (.I(net672),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output673 (.I(net673),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output674 (.I(net674),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output675 (.I(net675),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout676 (.I(net677),
    .Z(net676));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout677 (.I(net680),
    .Z(net677));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout678 (.I(net679),
    .Z(net678));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout679 (.I(net680),
    .Z(net679));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout680 (.I(net684),
    .Z(net680));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout681 (.I(net683),
    .Z(net681));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout682 (.I(net683),
    .Z(net682));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout683 (.I(net684),
    .Z(net683));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout684 (.I(net685),
    .Z(net684));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout685 (.I(net686),
    .Z(net685));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout686 (.I(net415),
    .Z(net686));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout687 (.I(net688),
    .Z(net687));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout688 (.I(net689),
    .Z(net688));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout689 (.I(net690),
    .Z(net689));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout690 (.I(net473),
    .Z(net690));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout691 (.I(net693),
    .Z(net691));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout692 (.I(net693),
    .Z(net692));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout693 (.I(net440),
    .Z(net693));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout694 (.I(net53),
    .Z(net694));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout695 (.I(net46),
    .Z(net695));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout696 (.I(net45),
    .Z(net696));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout697 (.I(net44),
    .Z(net697));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout698 (.I(net43),
    .Z(net698));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout699 (.I(net42),
    .Z(net699));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout700 (.I(net702),
    .Z(net700));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout701 (.I(net702),
    .Z(net701));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout702 (.I(net704),
    .Z(net702));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout703 (.I(net704),
    .Z(net703));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout704 (.I(net705),
    .Z(net704));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout705 (.I(net706),
    .Z(net705));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout706 (.I(net710),
    .Z(net706));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout707 (.I(net709),
    .Z(net707));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout708 (.I(net709),
    .Z(net708));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout709 (.I(net710),
    .Z(net709));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout710 (.I(net711),
    .Z(net710));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout711 (.I(net343),
    .Z(net711));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_712 (.ZN(net712));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0882__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0873__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0864__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0928__I (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0919__I (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0910__I (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0901__I (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__S (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0933__S (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0931__S (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0929__S (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0966__I (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0956__I (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0947__I (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0938__I (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0964__S (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__S (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0959__S (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__S (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0962__I (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0965__I (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0973__S (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0971__S (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0969__S (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__S (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0968__I (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1010__I (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0988__I (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0984__I (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0983__I (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0994__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0990__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0986__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1026__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1018__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1009__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__A2 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__A2 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0997__A2 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0993__A2 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A2 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1015__A3 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1006__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__A2 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1000__A2 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1025__A2 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1020__S (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1017__A2 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1002__S (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1036__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1032__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1028__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1037__A1 (.I(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1033__A1 (.I(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1029__A1 (.I(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__A1 (.I(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__A3 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__A1 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1016__I (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1030__A2 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1022__A2 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1019__A2 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1018__A3 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1058__I (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1054__I (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1040__I (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1039__I (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1053__A1 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1049__A1 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1045__A1 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1042__A2 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1048__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1044__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1041__A2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1071__A1 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1067__A1 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1063__A1 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1060__A1 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__A2 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1056__A2 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1070__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1066__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1062__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1059__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1041__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0924__I0 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0448__I0 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0920__I0 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0458__S0 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0451__S0 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0445__S0 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1038__A2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0922__I0 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0451__S1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0445__S1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0464__S (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0459__S (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0452__S (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0448__S (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1044__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0926__I0 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0452__I0 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1048__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0993__A1 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0929__I0 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0459__I0 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__A3 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1047__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0533__I0 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0458__I2 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0995__A3 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0992__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0555__I0 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0458__I3 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0473__S1 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0468__S1 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0463__S1 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0458__S1 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0997__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0931__I0 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0464__I0 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0478__S0 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0473__S0 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0468__S0 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0463__S0 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1059__A1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1002__I1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0933__I0 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0470__I0 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1000__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0559__I0 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0468__I3 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0483__S (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0479__S (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0474__S (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0470__S (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1062__A1 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__A1 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__I0 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0474__I0 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1066__A1 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__A1 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0939__I0 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0479__I0 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1014__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1011__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0564__I0 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0478__I3 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1070__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1017__A1 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__I0 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0483__I0 (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0917__I0 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0503__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0500__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0497__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0606__B1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0520__A2 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0517__A2 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0514__A2 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0520__B1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0517__B1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0514__B1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1046__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1043__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1042__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0526__I0 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0603__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0601__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0529__S (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0526__S (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1046__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1043__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0529__I0 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0590__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0581__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0568__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0532__I (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0540__S (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0537__S (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0535__S (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0533__S (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1068__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1064__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1061__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0540__I0 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0552__S (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0549__S (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0546__S (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0544__S (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0991__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0987__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0986__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0549__I0 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0995__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0991__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0987__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0552__I0 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0609__S (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0607__S (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0566__S (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0564__S (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0570__I (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__S (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0640__S (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0638__S (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0575__I (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__I0 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0606__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0600__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0576__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1038__A3 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0981__A2 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__A2 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0606__B2 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0618__S (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0616__S (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0614__S (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0612__S (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0627__S (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0625__S (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0623__S (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0621__S (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0636__S (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0634__S (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0632__S (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0630__S (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0646__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0651__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0662__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0656__A4 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0662__A3 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0661__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0661__A4 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0662__A4 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0684__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0667__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0683__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0672__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0683__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0677__A3 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0677__A4 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0683__A3 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0682__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0682__A4 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0684__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0979__S (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0975__S (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0775__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0686__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0718__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0716__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0714__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0687__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__I (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0740__I (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0697__I (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0690__I (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0784__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0695__S (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0693__S (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0691__S (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0731__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0722__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0707__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0698__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0720__S (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0712__S (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0710__S (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0708__S (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0738__S (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0736__S (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0734__S (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0732__S (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0768__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0759__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0750__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0741__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0786__S (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0773__S (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0771__S (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0769__S (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0816__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0807__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0798__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0789__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0796__S (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0794__S (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0792__S (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0790__S (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0823__S (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0821__S (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0819__S (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0817__S (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0937__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0900__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0863__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0826__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0854__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0845__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0836__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0827__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1055__A1 (.I(\data_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__A1 (.I(\data_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0523__I (.I(\data_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0445__I2 (.I(\data_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1055__A2 (.I(\data_load_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0528__I (.I(\data_load_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0451__I2 (.I(\data_load_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1055__A4 (.I(\data_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1051__A1 (.I(\data_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0535__I0 (.I(\data_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0463__I2 (.I(\data_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__A1 (.I(\data_load_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1056__A1 (.I(\data_load_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0537__I0 (.I(\data_load_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0468__I2 (.I(\data_load_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1069__A1 (.I(\data_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0546__I0 (.I(\data_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0482__I2 (.I(\data_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(data_read_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(data_read_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(data_read_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(data_read_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(data_read_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(data_read_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(data_read_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(data_read_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(data_read_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(data_read_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(data_read_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(data_read_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(data_read_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(data_read_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(data_read_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(data_read_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(hlt));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(instr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(instr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(instr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(instr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(instr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(instr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(instr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(instr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(instr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(instr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(instr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(instr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(instr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(instr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(instr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(instr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0999__A1 (.I(\instr_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0995__A1 (.I(\instr_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0548__I (.I(\instr_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0445__I3 (.I(\instr_load_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__A1 (.I(\instr_load_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1030__A1 (.I(\instr_load_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1027__A1 (.I(\instr_load_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0501__A1 (.I(\instr_load_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__A2 (.I(\instr_load_addr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1031__A1 (.I(\instr_load_addr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0505__A1 (.I(\instr_load_addr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1035__A1 (.I(\instr_load_addr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0509__A1 (.I(\instr_load_addr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0999__A2 (.I(\instr_load_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0551__I (.I(\instr_load_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0451__I3 (.I(\instr_load_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0999__A4 (.I(\instr_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0996__A1 (.I(\instr_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0557__I0 (.I(\instr_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0463__I3 (.I(\instr_load_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__A2 (.I(\instr_load_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__B (.I(\instr_load_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0561__I0 (.I(\instr_load_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0473__I3 (.I(\instr_load_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1015__A2 (.I(\instr_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1014__B (.I(\instr_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0566__I0 (.I(\instr_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0482__I3 (.I(\instr_load_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(io_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(io_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(io_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(io_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(io_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(io_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(io_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(io_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(io_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(io_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(io_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(io_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(io_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(io_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(io_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(io_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(la_data_in[100]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(la_data_in[101]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(la_data_in[102]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(la_data_in[103]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(la_data_in[104]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(la_data_in[105]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(la_data_in[106]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(la_data_in[107]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(la_data_in[108]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(la_data_in[109]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(la_data_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(la_data_in[110]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(la_data_in[111]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(la_data_in[112]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(la_data_in[113]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(la_data_in[114]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(la_data_in[115]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(la_data_in[116]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(la_data_in[117]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(la_data_in[118]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(la_data_in[119]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(la_data_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(la_data_in[120]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(la_data_in[121]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(la_data_in[122]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(la_data_in[123]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(la_data_in[124]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(la_data_in[125]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(la_data_in[126]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(la_data_in[127]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(la_data_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(la_data_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(la_data_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(la_data_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(la_data_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(la_data_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(la_data_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(la_data_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(la_data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(la_data_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input95_I (.I(la_data_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(la_data_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(la_data_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input98_I (.I(la_data_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input99_I (.I(la_data_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input100_I (.I(la_data_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input101_I (.I(la_data_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input102_I (.I(la_data_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input103_I (.I(la_data_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input104_I (.I(la_data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input105_I (.I(la_data_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input106_I (.I(la_data_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input107_I (.I(la_data_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input108_I (.I(la_data_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input109_I (.I(la_data_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input110_I (.I(la_data_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input111_I (.I(la_data_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input112_I (.I(la_data_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input113_I (.I(la_data_in[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input114_I (.I(la_data_in[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input115_I (.I(la_data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input116_I (.I(la_data_in[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input117_I (.I(la_data_in[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input118_I (.I(la_data_in[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input119_I (.I(la_data_in[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input120_I (.I(la_data_in[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input121_I (.I(la_data_in[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input122_I (.I(la_data_in[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input123_I (.I(la_data_in[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input124_I (.I(la_data_in[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input125_I (.I(la_data_in[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input126_I (.I(la_data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input127_I (.I(la_data_in[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input128_I (.I(la_data_in[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input129_I (.I(la_data_in[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input130_I (.I(la_data_in[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input131_I (.I(la_data_in[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input132_I (.I(la_data_in[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input133_I (.I(la_data_in[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input134_I (.I(la_data_in[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input135_I (.I(la_data_in[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input136_I (.I(la_data_in[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input137_I (.I(la_data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input138_I (.I(la_data_in[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input139_I (.I(la_data_in[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input140_I (.I(la_data_in[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input141_I (.I(la_data_in[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input142_I (.I(la_data_in[64]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input143_I (.I(la_data_in[65]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input144_I (.I(la_data_in[66]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input145_I (.I(la_data_in[67]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input146_I (.I(la_data_in[68]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input147_I (.I(la_data_in[69]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input148_I (.I(la_data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input149_I (.I(la_data_in[70]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input150_I (.I(la_data_in[71]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input151_I (.I(la_data_in[72]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input152_I (.I(la_data_in[73]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input153_I (.I(la_data_in[74]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input154_I (.I(la_data_in[75]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input155_I (.I(la_data_in[76]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input156_I (.I(la_data_in[77]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input157_I (.I(la_data_in[78]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input158_I (.I(la_data_in[79]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input159_I (.I(la_data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input160_I (.I(la_data_in[80]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input161_I (.I(la_data_in[81]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input162_I (.I(la_data_in[82]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input163_I (.I(la_data_in[83]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input164_I (.I(la_data_in[84]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input165_I (.I(la_data_in[85]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input166_I (.I(la_data_in[86]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input167_I (.I(la_data_in[87]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input168_I (.I(la_data_in[88]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input169_I (.I(la_data_in[89]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input170_I (.I(la_data_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input171_I (.I(la_data_in[90]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input172_I (.I(la_data_in[91]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input173_I (.I(la_data_in[92]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input174_I (.I(la_data_in[93]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input175_I (.I(la_data_in[94]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input176_I (.I(la_data_in[95]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input177_I (.I(la_data_in[96]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input178_I (.I(la_data_in[97]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input179_I (.I(la_data_in[98]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input180_I (.I(la_data_in[99]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input181_I (.I(la_data_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input182_I (.I(la_oenb[100]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input183_I (.I(la_oenb[101]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input184_I (.I(la_oenb[102]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input185_I (.I(la_oenb[103]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input186_I (.I(la_oenb[104]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input187_I (.I(la_oenb[105]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input188_I (.I(la_oenb[106]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input189_I (.I(la_oenb[107]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input190_I (.I(la_oenb[108]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input191_I (.I(la_oenb[109]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input192_I (.I(la_oenb[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input193_I (.I(la_oenb[110]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input194_I (.I(la_oenb[111]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input195_I (.I(la_oenb[112]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input196_I (.I(la_oenb[113]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input197_I (.I(la_oenb[114]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input198_I (.I(la_oenb[115]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input199_I (.I(la_oenb[116]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input200_I (.I(la_oenb[117]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input201_I (.I(la_oenb[118]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input202_I (.I(la_oenb[119]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input203_I (.I(la_oenb[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input204_I (.I(la_oenb[120]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input205_I (.I(la_oenb[121]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input206_I (.I(la_oenb[122]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input207_I (.I(la_oenb[123]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input208_I (.I(la_oenb[124]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input209_I (.I(la_oenb[125]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input210_I (.I(la_oenb[126]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input211_I (.I(la_oenb[127]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input212_I (.I(la_oenb[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input213_I (.I(la_oenb[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input214_I (.I(la_oenb[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input215_I (.I(la_oenb[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input216_I (.I(la_oenb[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input217_I (.I(la_oenb[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input218_I (.I(la_oenb[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input219_I (.I(la_oenb[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input220_I (.I(la_oenb[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input221_I (.I(la_oenb[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input222_I (.I(la_oenb[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input223_I (.I(la_oenb[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input224_I (.I(la_oenb[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input225_I (.I(la_oenb[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input226_I (.I(la_oenb[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input227_I (.I(la_oenb[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input228_I (.I(la_oenb[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input229_I (.I(la_oenb[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input230_I (.I(la_oenb[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input231_I (.I(la_oenb[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input232_I (.I(la_oenb[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input233_I (.I(la_oenb[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input234_I (.I(la_oenb[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input235_I (.I(la_oenb[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input236_I (.I(la_oenb[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input237_I (.I(la_oenb[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input238_I (.I(la_oenb[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input239_I (.I(la_oenb[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input240_I (.I(la_oenb[38]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input241_I (.I(la_oenb[39]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input242_I (.I(la_oenb[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input243_I (.I(la_oenb[40]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input244_I (.I(la_oenb[41]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input245_I (.I(la_oenb[42]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input246_I (.I(la_oenb[43]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input247_I (.I(la_oenb[44]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input248_I (.I(la_oenb[45]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input249_I (.I(la_oenb[46]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input250_I (.I(la_oenb[47]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input251_I (.I(la_oenb[48]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input252_I (.I(la_oenb[49]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input253_I (.I(la_oenb[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input254_I (.I(la_oenb[50]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input255_I (.I(la_oenb[51]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input256_I (.I(la_oenb[52]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input257_I (.I(la_oenb[53]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input258_I (.I(la_oenb[54]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input259_I (.I(la_oenb[55]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input260_I (.I(la_oenb[56]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input261_I (.I(la_oenb[57]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input262_I (.I(la_oenb[58]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input263_I (.I(la_oenb[59]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input264_I (.I(la_oenb[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input265_I (.I(la_oenb[60]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input266_I (.I(la_oenb[61]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input267_I (.I(la_oenb[62]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input268_I (.I(la_oenb[63]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input269_I (.I(la_oenb[64]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input270_I (.I(la_oenb[65]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input271_I (.I(la_oenb[66]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input272_I (.I(la_oenb[67]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input273_I (.I(la_oenb[68]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input274_I (.I(la_oenb[69]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input275_I (.I(la_oenb[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input276_I (.I(la_oenb[70]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input277_I (.I(la_oenb[71]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input278_I (.I(la_oenb[72]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input279_I (.I(la_oenb[73]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input280_I (.I(la_oenb[74]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input281_I (.I(la_oenb[75]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input282_I (.I(la_oenb[76]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input283_I (.I(la_oenb[77]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input284_I (.I(la_oenb[78]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input285_I (.I(la_oenb[79]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input286_I (.I(la_oenb[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input287_I (.I(la_oenb[80]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input288_I (.I(la_oenb[81]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input289_I (.I(la_oenb[82]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input290_I (.I(la_oenb[83]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input291_I (.I(la_oenb[84]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input292_I (.I(la_oenb[85]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input293_I (.I(la_oenb[86]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input294_I (.I(la_oenb[87]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input295_I (.I(la_oenb[88]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input296_I (.I(la_oenb[89]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input297_I (.I(la_oenb[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input298_I (.I(la_oenb[90]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input299_I (.I(la_oenb[91]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input300_I (.I(la_oenb[92]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input301_I (.I(la_oenb[93]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input302_I (.I(la_oenb[94]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input303_I (.I(la_oenb[95]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input304_I (.I(la_oenb[96]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input305_I (.I(la_oenb[97]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input306_I (.I(la_oenb[98]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input307_I (.I(la_oenb[99]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input308_I (.I(la_oenb[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input309_I (.I(uP_data_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input310_I (.I(uP_data_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input311_I (.I(uP_data_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input312_I (.I(uP_data_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input313_I (.I(uP_data_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input314_I (.I(uP_data_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input315_I (.I(uP_data_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input316_I (.I(uP_data_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input317_I (.I(uP_dataw_en));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input318_I (.I(uP_instr_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input319_I (.I(uP_instr_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input320_I (.I(uP_instr_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input321_I (.I(uP_instr_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input322_I (.I(uP_instr_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input323_I (.I(uP_instr_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input324_I (.I(uP_instr_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input325_I (.I(uP_instr_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input326_I (.I(uP_write_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input327_I (.I(uP_write_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input328_I (.I(uP_write_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input329_I (.I(uP_write_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input330_I (.I(uP_write_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input331_I (.I(uP_write_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input332_I (.I(uP_write_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input333_I (.I(uP_write_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input334_I (.I(uP_write_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input335_I (.I(uP_write_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input336_I (.I(uP_write_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input337_I (.I(uP_write_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input338_I (.I(uP_write_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input339_I (.I(uP_write_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input340_I (.I(uP_write_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input341_I (.I(uP_write_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input342_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input343_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input344_I (.I(wbs_adr_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input345_I (.I(wbs_adr_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input346_I (.I(wbs_adr_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input347_I (.I(wbs_adr_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input348_I (.I(wbs_adr_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input349_I (.I(wbs_adr_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input350_I (.I(wbs_adr_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input351_I (.I(wbs_adr_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input352_I (.I(wbs_adr_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input353_I (.I(wbs_adr_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input354_I (.I(wbs_adr_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input355_I (.I(wbs_adr_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input356_I (.I(wbs_adr_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input357_I (.I(wbs_adr_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input358_I (.I(wbs_adr_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input359_I (.I(wbs_adr_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input360_I (.I(wbs_adr_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input361_I (.I(wbs_adr_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input362_I (.I(wbs_adr_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input363_I (.I(wbs_adr_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input364_I (.I(wbs_adr_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input365_I (.I(wbs_adr_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input366_I (.I(wbs_adr_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input367_I (.I(wbs_adr_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input368_I (.I(wbs_adr_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input369_I (.I(wbs_adr_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input370_I (.I(wbs_adr_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input371_I (.I(wbs_adr_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input372_I (.I(wbs_adr_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input373_I (.I(wbs_adr_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input374_I (.I(wbs_adr_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input375_I (.I(wbs_adr_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input376_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input377_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input378_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input379_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input380_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input381_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input382_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input383_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input384_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input385_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input386_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input387_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input388_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input389_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input390_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input391_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input392_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input393_I (.I(wbs_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input394_I (.I(wbs_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input395_I (.I(wbs_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input396_I (.I(wbs_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input397_I (.I(wbs_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input398_I (.I(wbs_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input399_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input400_I (.I(wbs_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input401_I (.I(wbs_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input402_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input403_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input404_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input405_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input406_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input407_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input408_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input409_I (.I(wbs_sel_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input410_I (.I(wbs_sel_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input411_I (.I(wbs_sel_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input412_I (.I(wbs_sel_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input413_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input414_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0823__I0 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0445__I0 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0848__I0 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0501__B2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0850__I0 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0505__B2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0852__I0 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0509__B2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0855__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0514__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0857__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0517__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0859__I0 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0520__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0828__I0 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0451__I0 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0830__I0 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0458__I0 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0832__I0 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0463__I0 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0834__I0 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0468__I0 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0837__I0 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0473__I0 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0839__I0 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0478__I0 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0841__I0 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0482__I0 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0843__I0 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0494__B2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0846__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0498__B2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0569__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0445__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0593__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0501__C2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0595__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0505__C2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0597__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0509__C2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0599__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0514__B2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0601__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0517__B2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0603__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0520__B2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0571__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0451__I1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0573__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0458__I1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0577__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0463__I1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0579__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0468__I1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0582__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0473__I1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0584__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0478__I1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0586__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0482__I1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0588__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0494__C2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0591__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0498__C2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1199__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0607__I0 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0440__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1200__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0609__I0 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0450__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1201__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0612__I0 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0454__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1202__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0614__I0 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0461__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1203__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0616__I0 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0466__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1204__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0618__I0 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0472__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1205__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0621__I0 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0476__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1206__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0623__I0 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0481__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout699_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout698_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1208__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout697_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout696_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1210__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout695_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0954__I0 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0636__I0 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0515__A2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__I0 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0638__I0 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0518__A2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1214__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0959__I0 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0640__I0 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0521__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0495__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0485__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0446__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0491__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0489__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0441__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0492__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0489__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0457__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0443__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout694_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1225__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__I0 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0973__I0 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__I1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0964__I1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__I1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0526__I1 (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0529__I1 (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0533__I1 (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0535__I1 (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0537__I1 (.I(net313));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0540__I1 (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0544__I1 (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0546__I1 (.I(net316));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0969__I0 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0606__A2 (.I(net317));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0549__I1 (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0552__I1 (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0555__I1 (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0557__I1 (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__I1 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0975__I0 (.I(net342));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout711_I (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__I (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__I (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1173__I (.I(net346));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1174__I (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1175__I (.I(net348));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1176__I (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1177__I (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__I (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1179__I (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1180__I (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1181__I (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1163__I (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1183__I (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1184__I (.I(net358));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1185__I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__I (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1187__I (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1188__I (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__I (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1190__I (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0708__I0 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1164__I (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0710__I0 (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0712__I0 (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__I (.I(net369));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1166__I (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1167__I (.I(net371));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1168__I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1169__I (.I(net373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__I (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1171__I (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0703__I0 (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0691__I0 (.I(net409));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0693__I0 (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0695__I0 (.I(net411));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0699__I0 (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0705__I0 (.I(net413));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0701__I0 (.I(net414));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output416_I (.I(net416));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0861__I0 (.I(net416));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output417_I (.I(net417));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0865__I0 (.I(net417));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output418_I (.I(net418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0867__I0 (.I(net418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output419_I (.I(net419));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0869__I0 (.I(net419));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output420_I (.I(net420));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0871__I0 (.I(net420));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output421_I (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0874__I0 (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output422_I (.I(net422));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0876__I0 (.I(net422));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output423_I (.I(net423));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0878__I0 (.I(net423));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output424_I (.I(net424));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0786__I0 (.I(net424));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output425_I (.I(net425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0810__I0 (.I(net425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output426_I (.I(net426));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0812__I0 (.I(net426));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output427_I (.I(net427));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0814__I0 (.I(net427));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output428_I (.I(net428));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0817__I0 (.I(net428));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output429_I (.I(net429));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0819__I0 (.I(net429));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output430_I (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0821__I0 (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output431_I (.I(net431));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0790__I0 (.I(net431));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output432_I (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0792__I0 (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output433_I (.I(net433));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0794__I0 (.I(net433));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output434_I (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0796__I0 (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output435_I (.I(net435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0799__I0 (.I(net435));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output436_I (.I(net436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0801__I0 (.I(net436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output437_I (.I(net437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0803__I0 (.I(net437));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output438_I (.I(net438));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0805__I0 (.I(net438));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output439_I (.I(net439));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0808__I0 (.I(net439));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout693_I (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1198__I (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output449_I (.I(net449));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0757__I0 (.I(net449));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output450_I (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0760__I0 (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output451_I (.I(net451));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0762__I0 (.I(net451));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output452_I (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0764__I0 (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output453_I (.I(net453));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0766__I0 (.I(net453));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output454_I (.I(net454));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0769__I0 (.I(net454));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output455_I (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0771__I0 (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output456_I (.I(net456));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0773__I0 (.I(net456));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output460_I (.I(net460));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output461_I (.I(net461));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output462_I (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output463_I (.I(net463));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output464_I (.I(net464));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output467_I (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output468_I (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output469_I (.I(net469));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output470_I (.I(net470));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output480_I (.I(net480));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output481_I (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output482_I (.I(net482));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0880__I0 (.I(net482));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output483_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0904__I0 (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output484_I (.I(net484));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0906__I0 (.I(net484));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output485_I (.I(net485));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0908__I0 (.I(net485));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output486_I (.I(net486));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0911__I0 (.I(net486));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output487_I (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0913__I0 (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output488_I (.I(net488));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0915__I0 (.I(net488));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output489_I (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0883__I0 (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output490_I (.I(net490));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0885__I0 (.I(net490));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output491_I (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output492_I (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0887__I0 (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output493_I (.I(net493));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0889__I0 (.I(net493));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output494_I (.I(net494));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0892__I0 (.I(net494));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output495_I (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__I0 (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output496_I (.I(net496));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0896__I0 (.I(net496));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output497_I (.I(net497));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0898__I0 (.I(net497));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output498_I (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0902__I0 (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output521_I (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output522_I (.I(net522));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output625_I (.I(net625));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output626_I (.I(net626));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output627_I (.I(net627));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0720__I0 (.I(net627));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output628_I (.I(net628));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0744__I0 (.I(net628));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output629_I (.I(net629));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0746__I0 (.I(net629));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output630_I (.I(net630));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0748__I0 (.I(net630));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output631_I (.I(net631));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0751__I0 (.I(net631));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output632_I (.I(net632));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0753__I0 (.I(net632));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output633_I (.I(net633));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0755__I0 (.I(net633));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output634_I (.I(net634));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0723__I0 (.I(net634));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output635_I (.I(net635));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0725__I0 (.I(net635));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output636_I (.I(net636));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0727__I0 (.I(net636));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output637_I (.I(net637));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0729__I0 (.I(net637));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output638_I (.I(net638));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0732__I0 (.I(net638));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output639_I (.I(net639));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0734__I0 (.I(net639));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output640_I (.I(net640));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0736__I0 (.I(net640));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output641_I (.I(net641));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0738__I0 (.I(net641));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output642_I (.I(net642));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0742__I0 (.I(net642));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output643_I (.I(net643));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1090__CLK (.I(net677));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1077__CLK (.I(net677));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1089__CLK (.I(net677));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout676_I (.I(net677));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout679_I (.I(net680));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout677_I (.I(net680));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1082__CLK (.I(net681));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1081__CLK (.I(net681));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1093__CLK (.I(net681));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1080__CLK (.I(net681));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout683_I (.I(net684));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout680_I (.I(net684));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1086__CLK (.I(net685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1085__CLK (.I(net685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1084__CLK (.I(net685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout684_I (.I(net685));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout685_I (.I(net686));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output415_I (.I(net686));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0979__I0 (.I(net686));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout689_I (.I(net690));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output473_I (.I(net690));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__I (.I(net690));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1215__I (.I(net690));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output440_I (.I(net691));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1193__I (.I(net691));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1192__I (.I(net691));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__I (.I(net691));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1196__I (.I(net692));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1195__I (.I(net692));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1194__I (.I(net692));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1197__I (.I(net693));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__I0 (.I(net693));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout691_I (.I(net693));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout692_I (.I(net693));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0605__A2 (.I(net694));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0524__I (.I(net694));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0542__I (.I(net694));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0531__I (.I(net694));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1036__A1 (.I(net695));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0634__I0 (.I(net695));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0510__A2 (.I(net695));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0952__I0 (.I(net695));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1032__A1 (.I(net696));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0632__I0 (.I(net696));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0507__A2 (.I(net696));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0950__I0 (.I(net696));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1028__A1 (.I(net697));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0630__I0 (.I(net697));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0502__A2 (.I(net697));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0948__I0 (.I(net697));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1025__A1 (.I(net698));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0627__I0 (.I(net698));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0499__A2 (.I(net698));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0945__I0 (.I(net698));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1020__I1 (.I(net699));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0625__I0 (.I(net699));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0496__A2 (.I(net699));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0943__I0 (.I(net699));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1079__RN (.I(net702));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1074__RN (.I(net702));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout700_I (.I(net702));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout701_I (.I(net702));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout702_I (.I(net704));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout703_I (.I(net704));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1092__RN (.I(net705));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1080__RN (.I(net705));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1078__RN (.I(net705));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout704_I (.I(net705));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1093__RN (.I(net706));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout705_I (.I(net706));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1094__RN (.I(net707));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1083__RN (.I(net707));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1082__RN (.I(net707));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1081__RN (.I(net707));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout707_I (.I(net709));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout708_I (.I(net709));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout709_I (.I(net710));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout706_I (.I(net710));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout710_I (.I(net711));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1224__I (.I(net711));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0971__I0 (.I(net711));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3187 ();
 assign Serial_output = net712;
 assign data_mem_sel = net713;
 assign instr_mem_sel = net714;
 assign io_oeb[0] = net715;
 assign io_oeb[10] = net725;
 assign io_oeb[11] = net726;
 assign io_oeb[12] = net727;
 assign io_oeb[13] = net728;
 assign io_oeb[14] = net729;
 assign io_oeb[15] = net730;
 assign io_oeb[16] = net758;
 assign io_oeb[17] = net759;
 assign io_oeb[18] = net760;
 assign io_oeb[19] = net761;
 assign io_oeb[1] = net716;
 assign io_oeb[20] = net762;
 assign io_oeb[21] = net763;
 assign io_oeb[22] = net764;
 assign io_oeb[23] = net765;
 assign io_oeb[24] = net766;
 assign io_oeb[25] = net767;
 assign io_oeb[26] = net768;
 assign io_oeb[27] = net769;
 assign io_oeb[28] = net770;
 assign io_oeb[29] = net771;
 assign io_oeb[2] = net717;
 assign io_oeb[30] = net772;
 assign io_oeb[31] = net773;
 assign io_oeb[32] = net774;
 assign io_oeb[33] = net775;
 assign io_oeb[34] = net776;
 assign io_oeb[35] = net731;
 assign io_oeb[36] = net777;
 assign io_oeb[37] = net778;
 assign io_oeb[3] = net718;
 assign io_oeb[4] = net719;
 assign io_oeb[5] = net720;
 assign io_oeb[6] = net721;
 assign io_oeb[7] = net722;
 assign io_oeb[8] = net723;
 assign io_oeb[9] = net724;
 assign io_out[16] = net732;
 assign io_out[17] = net733;
 assign io_out[18] = net734;
 assign io_out[19] = net735;
 assign io_out[20] = net736;
 assign io_out[21] = net737;
 assign io_out[22] = net738;
 assign io_out[23] = net739;
 assign io_out[24] = net740;
 assign io_out[25] = net741;
 assign io_out[26] = net742;
 assign io_out[27] = net743;
 assign io_out[28] = net744;
 assign io_out[29] = net745;
 assign io_out[30] = net746;
 assign io_out[31] = net747;
 assign io_out[32] = net748;
 assign io_out[33] = net749;
 assign io_out[34] = net750;
 assign io_out[36] = net751;
 assign io_out[37] = net752;
 assign irq[0] = net753;
 assign irq[1] = net754;
 assign irq[2] = net755;
 assign la_data_out[0] = net756;
 assign la_data_out[1] = net757;
endmodule

